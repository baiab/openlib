
.subckt BUFTD1  I OE Z
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.14175p as=0.1053p l=0.09u nrd=0.702 nrs=0.52 pd=1.854u ps=1.368u sa=2.115e-07 sb=2.34e-07 w=0.45u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.03726p as=0.03159p l=0.09u nrd=0.509 nrs=0.433 pd=0.693u ps=0.504u sa=4.86e-07 sb=7.695e-07 w=0.27u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.08991p as=0.0324p l=0.09u nrd=0.696 nrs=0.25 pd=1.1313u ps=0.54u sa=3.465e-07 sb=4.77e-07 w=0.36u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.07452p as=0.0324p l=0.09u nrd=0.575 nrs=0.25 pd=1.134u ps=0.54u sa=6.795e-07 sb=2.07e-07 w=0.36u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.05589p as=0.03726p l=0.09u nrd=0.767 nrs=0.509 pd=0.954u ps=0.693u sa=2.07e-07 sb=1.0737e-06 w=0.27u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.03159p as=0.06804p l=0.09u nrd=0.433 nrs=0.929 pd=0.504u ps=0.8487u sa=8.1e-07 sb=3.834e-07 w=0.27u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK pch ad=0.07452p as=0.06723p l=0.09u nrd=0.575 nrs=0.52 pd=1.134u ps=0.828u sa=2.07e-07 sb=7.83e-07 w=0.36u 
MM9 M9:DRN M9:GATE M9:SRC M9:BULK pch ad=0.0648p as=0.14904p l=0.09u nrd=0.125 nrs=0.287 pd=0.9u ps=1.854u sa=5.985e-07 sb=2.07e-07 w=0.72u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK pch ad=0.10692p as=0.04212p l=0.09u nrd=0.822 nrs=0.325 pd=1.53u ps=0.594u sa=2.07e-07 sb=8.91e-07 w=0.36u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK pch ad=0.12312p as=0.13041p l=0.09u nrd=0.31 nrs=0.329 pd=1.3977u ps=1.674u sa=4.104e-07 sb=2.07e-07 w=0.63u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK pch ad=0.13446p as=0.0648p l=0.09u nrd=0.26 nrs=0.125 pd=1.656u ps=0.9u sa=3.015e-07 sb=4.77e-07 w=0.72u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK pch ad=0.04212p as=0.07047p l=0.09u nrd=0.325 nrs=0.543 pd=0.594u ps=0.7983u sa=5.31e-07 sb=5.67e-07 w=0.36u 
R1 M6:BULK M4:DRN 2.18524e-05
R2 M6:BULK M3:BULK 0.001
R3 M6:BULK M4:BULK 0.001
R4 M6:BULK M5:BULK 0.001
R5 M6:BULK M1:BULK 0.001
R6 M6:BULK M2:BULK 0.001
R7 M5:SRC M6:DRN 2.27273e-10
R8 M5:SRC M4:DRN 6.72554e-10
R9 M4:DRN GND 1.64127
R10 M4:DRN M3:SRC 0.001
R11 M4:DRN M2:DRN 0.001
R12 M12:SRC Z 9.34108
R13 Z M2:SRC 18.2965
R14 M12:GATE M1:DRN 158.763
R15 M12:GATE M11:DRN 159.275
R16 M11:DRN M1:DRN 41.9253
R17 M11:DRN M10:SRC 0.001
R18 M9:SRC M5:DRN 43.127
R19 M9:SRC M2:GATE 130.5
R20 M2:GATE M5:DRN 124.958
R21 M5:DRN M4:SRC 0.001
R22 M11:GATE OE 162.614
R23 M11:GATE M1:GATE 358.174
R24 M7:GATE M3:GATE 245.258
R25 M7:GATE OE 57.1884
R26 OE M3:GATE 109.838
R27 OE M1:GATE 58.409
R28 M1:SRC M6:SRC 0.001
R29 M8:GATE M3:DRN 406.639
R30 M8:GATE M4:GATE 230.459
R31 M8:GATE M7:DRN 413.273
R32 M7:DRN M3:DRN 45.8192
R33 M7:DRN M4:GATE 118.951
R34 M3:DRN M4:GATE 117.041
R35 M9:DRN M8:SRC 0.001
R36 I:1 M5:GATE 63.6
R37 I:1 I 33.1975
R38 I:1 M6:GATE 79.9395
R39 I:1 M9:GATE 71.28
R40 I:1 M10:GATE 248.981
R41 M10:GATE I 317.827
R42 M10:GATE M6:GATE 765.326
R43 I M6:GATE 102.044
R44 M12:BULK M8:BULK 0.001
R45 M12:BULK M8:DRN 2.18516e-05
R46 M12:BULK M10:DRN 0.00342936
R47 M12:BULK M9:BULK 0.001
R48 M12:BULK M12:DRN 0.00308642
R49 M12:BULK M7:BULK 0.001
R50 M12:BULK M10:BULK 0.001
R51 M12:BULK M11:BULK 0.001
R52 M10:DRN VDD 6.68523
R53 M10:DRN M8:DRN 1.22222e-09
R54 M10:DRN M12:DRN 2.1e-09
R55 VDD M8:DRN 3.13592
R56 VDD M12:DRN 5.10572
R57 M12:DRN M8:DRN 196.878
R58 M12:DRN M11:SRC 0.001
R59 M8:DRN M7:SRC 1.49425e-10
c_1 M5:SRC 0 2.23473e-20 
c_2 M6:DRN 0 2.90077e-19 
c_3 M4:DRN 0 1.10993e-16 
c_4 GND 0 8.32778e-17 
c_5 M12:SRC M4:DRN 2.75385e-19 
c_6 M12:SRC 0 6.34486e-18 
c_7 Z GND 2.6451e-17 
c_8 Z M4:DRN 9.9344e-19 
c_9 Z M6:BULK 7.64481e-18 
c_10 Z 0 4.2878e-17 
c_11 M2:SRC M5:SRC 1.35663e-19 
c_12 M2:SRC M4:DRN 1.02088e-17 
c_13 M2:SRC GND 1.80871e-18 
c_14 M2:SRC 0 1.23832e-18 
c_15 M12:GATE Z 5.60382e-17 
c_16 M12:GATE M12:SRC 3.40758e-17 
c_17 M12:GATE 0 2.04079e-17 
c_18 M11:DRN M4:DRN 4.55764e-20 
c_19 M11:DRN Z 1.7276e-17 
c_20 M11:DRN M12:SRC 3.28594e-19 
c_21 M1:DRN GND 4.23649e-18 
c_22 M1:DRN M4:DRN 2.57291e-17 
c_23 M1:DRN M2:SRC 1.20206e-18 
c_24 M1:DRN Z 6.59701e-18 
c_25 M1:DRN M5:SRC 3.04422e-19 
c_26 M1:DRN M12:SRC 7.97372e-19 
c_27 M1:DRN M6:DRN 1.73622e-20 
c_28 M1:DRN 0 2.56266e-19 
c_29 M9:SRC M4:DRN 2.15969e-20 
c_30 M9:SRC M1:DRN 8.57072e-18 
c_31 M9:SRC M5:SRC 1.03951e-19 
c_32 M9:SRC M6:BULK 1.80625e-17 
c_33 M9:SRC M11:DRN 1.00433e-16 
c_34 M9:SRC M12:SRC 6.24141e-20 
c_35 M9:SRC M6:DRN 2.0366e-18 
c_36 M2:GATE GND 6.81365e-18 
c_37 M2:GATE M4:DRN 2.53673e-17 
c_38 M2:GATE M2:SRC 1.82982e-17 
c_39 M2:GATE Z 7.60325e-17 
c_40 M2:GATE M6:BULK 1.96962e-18 
c_41 M2:GATE M11:DRN 2.35668e-17 
c_42 M2:GATE M12:GATE 4.01592e-18 
c_43 M2:GATE 0 1.89631e-17 
c_44 M5:DRN GND 1.86852e-16 
c_45 M5:DRN M4:DRN 4.02888e-17 
c_46 M5:DRN M1:DRN 7.64737e-18 
c_47 M5:DRN M5:SRC 2.7478e-18 
c_48 M5:DRN 0 3.71129e-19 
c_49 M11:GATE M4:DRN 1.76175e-19 
c_50 M11:GATE M2:GATE 4.01028e-18 
c_51 M11:GATE M9:SRC 7.97163e-19 
c_52 M11:GATE M11:DRN 3.98222e-17 
c_53 M11:GATE M12:GATE 3.93845e-18 
c_54 M11:GATE 0 1.19048e-17 
c_55 M7:GATE M5:DRN 1.33738e-18 
c_56 M7:GATE M6:BULK 5.34531e-18 
c_57 M7:GATE 0 1.6281e-18 
c_58 OE GND 1.1692e-18 
c_59 OE M4:DRN 2.85516e-18 
c_60 OE M5:DRN 4.02688e-20 
c_61 OE M1:DRN 1.68618e-16 
c_62 OE M9:SRC 1.15235e-16 
c_63 OE M6:BULK 1.99964e-17 
c_64 OE M11:DRN 4.0214e-18 
c_65 OE M12:GATE 2.72582e-18 
c_66 OE 0 2.10378e-18 
c_67 M1:GATE GND 2.72836e-18 
c_68 M1:GATE M4:DRN 8.47618e-18 
c_69 M1:GATE M1:DRN 1.40764e-17 
c_70 M1:GATE M2:GATE 1.14671e-20 
c_71 M1:GATE M9:SRC 2.03464e-17 
c_72 M1:GATE M5:SRC 5.66882e-19 
c_73 M1:GATE M6:BULK 1.19623e-18 
c_74 M1:GATE 0 7.65e-20 
c_75 M3:GATE M6:BULK 7.73228e-18 
c_76 M3:GATE M4:DRN 1.8202e-17 
c_77 M3:GATE M5:DRN 3.52247e-19 
c_78 M3:GATE GND 4.8844e-18 
c_79 M3:GATE 0 7.31108e-18 
c_80 M1:SRC M4:DRN 8.70522e-18 
c_81 M1:SRC M5:DRN 1.16999e-18 
c_82 M1:SRC GND 1.26933e-20 
c_83 M8:GATE M4:DRN 9.50298e-23 
c_84 M8:GATE OE 1.97901e-17 
c_85 M8:GATE M5:DRN 1.64733e-18 
c_86 M8:GATE M7:GATE 2.89756e-17 
c_87 M8:GATE M9:SRC 1.60689e-19 
c_88 M8:GATE 0 2.53956e-17 
c_89 M7:DRN OE 1.32158e-16 
c_90 M7:DRN M7:GATE 1.69539e-17 
c_91 M7:DRN M4:DRN 6.27184e-20 
c_92 M7:DRN 0 1.77695e-17 
c_93 M3:DRN GND 5.39816e-17 
c_94 M3:DRN M3:GATE 2.00676e-17 
c_95 M3:DRN M4:DRN 1.74722e-17 
c_96 M3:DRN M5:DRN 1.17048e-19 
c_97 M3:DRN M7:GATE 7.10557e-18 
c_98 M3:DRN M6:BULK 2.09335e-17 
c_99 M3:DRN M6:DRN 2.5472e-18 
c_100 M3:DRN 0 1.89498e-18 
c_101 M4:GATE GND 4.48678e-18 
c_102 M4:GATE M3:GATE 4.09845e-18 
c_103 M4:GATE M4:DRN 1.90284e-17 
c_104 M4:GATE M5:DRN 9.32231e-17 
c_105 M4:GATE M6:BULK 5.07854e-18 
c_106 M4:GATE M6:DRN 3.58477e-19 
c_107 M4:GATE 0 4.95758e-18 
c_108 M9:DRN OE 3.3296e-18 
c_109 M9:DRN M7:DRN 3.28594e-19 
c_110 M9:DRN M3:DRN 9.99708e-19 
c_111 M9:DRN M5:DRN 1.4291e-18 
c_112 I:1 GND 1.2173e-18 
c_113 I:1 M3:DRN 2.63202e-17 
c_114 I:1 M4:DRN 5.28241e-19 
c_115 I:1 M4:GATE 3.10712e-20 
c_116 I:1 OE 9.1877e-18 
c_117 I:1 M5:DRN 2.40831e-17 
c_118 I:1 M1:GATE 1.16215e-19 
c_119 I:1 M1:DRN 4.74511e-19 
c_120 I:1 M9:SRC 1.34693e-17 
c_121 I:1 M5:SRC 1.18568e-18 
c_122 I:1 M6:BULK 1.0032e-17 
c_123 I:1 M11:DRN 6.87378e-18 
c_124 I:1 M6:DRN 3.01681e-17 
c_125 M9:GATE OE 9.86544e-18 
c_126 M9:GATE M5:DRN 7.95584e-18 
c_127 M9:GATE M1:DRN 8.12522e-22 
c_128 M9:GATE M7:GATE 2.98035e-19 
c_129 M9:GATE M8:GATE 2.28085e-17 
c_130 M9:GATE M9:SRC 1.70591e-17 
c_131 M9:GATE M11:DRN 1.08584e-19 
c_132 M9:GATE M11:GATE 9.55943e-20 
c_133 M9:GATE 0 2.06949e-18 
c_134 M10:GATE M4:DRN 8.38719e-19 
c_135 M10:GATE OE 1.61293e-17 
c_136 M10:GATE M5:DRN 7.38947e-19 
c_137 M10:GATE M1:SRC 2.79941e-18 
c_138 M10:GATE M1:DRN 3.5242e-18 
c_139 M10:GATE M8:GATE 2.46895e-19 
c_140 M10:GATE M9:SRC 1.42256e-17 
c_141 M10:GATE M11:GATE 6.23273e-18 
c_142 M10:GATE M12:GATE 3.33686e-20 
c_143 M10:GATE 0 7.78539e-18 
c_144 I GND 1.58614e-18 
c_145 I M3:DRN 5.83791e-19 
c_146 I M4:DRN 1.54088e-18 
c_147 I OE 9.11442e-17 
c_148 I M1:DRN 1.50522e-17 
c_149 I M8:GATE 5.68677e-19 
c_150 I M9:SRC 7.99132e-17 
c_151 I M6:BULK 3.21005e-18 
c_152 I M11:DRN 1.09065e-17 
c_153 I 0 2.2897e-18 
c_154 M5:GATE M6:BULK 3.77171e-18 
c_155 M5:GATE M3:GATE 1.80529e-19 
c_156 M5:GATE M3:DRN 5.63023e-20 
c_157 M5:GATE M4:GATE 5.29967e-18 
c_158 M5:GATE M4:DRN 2.71009e-17 
c_159 M5:GATE M5:DRN 1.52278e-17 
c_160 M5:GATE GND 3.7055e-18 
c_161 M6:GATE GND 2.19511e-18 
c_162 M6:GATE M4:DRN 1.10998e-17 
c_163 M6:GATE M4:GATE 7.32822e-21 
c_164 M6:GATE OE 5.39935e-18 
c_165 M6:GATE M5:DRN 1.15087e-17 
c_166 M6:GATE M1:GATE 6.40137e-18 
c_167 M6:GATE M1:DRN 5.51652e-19 
c_168 M6:GATE M5:SRC 5.91843e-18 
c_169 M6:GATE M6:BULK 3.10788e-18 
c_170 M6:GATE M11:GATE 5.82797e-18 
c_171 M6:GATE 0 1.72161e-18 
c_172 M12:BULK M3:DRN 6.1463e-18 
c_173 M12:BULK M3:GATE 7.12986e-18 
c_174 M12:BULK OE 1.63451e-17 
c_175 M12:BULK I:1 7.23779e-18 
c_176 M12:BULK I 4.1277e-19 
c_177 M12:BULK M1:GATE 1.14283e-17 
c_178 M12:BULK Z 1.22532e-17 
c_179 M12:BULK M7:GATE 2.09951e-18 
c_180 M12:BULK M8:GATE 7.7976e-18 
c_181 M12:BULK M9:GATE 2.08394e-18 
c_182 M12:BULK M9:SRC 4.81448e-19 
c_183 M12:BULK M10:GATE 1.33927e-17 
c_184 M12:BULK M7:DRN 3.36069e-18 
c_185 M12:BULK M11:DRN 1.83161e-17 
c_186 M12:BULK M11:GATE 6.55169e-18 
c_187 M12:BULK M12:SRC 5.57072e-18 
c_188 M12:BULK M12:GATE 3.02274e-18 
c_189 M10:DRN OE 2.25972e-18 
c_190 M10:DRN I:1 7.8687e-18 
c_191 M10:DRN M1:DRN 4.91395e-19 
c_192 M10:DRN Z 8.10111e-20 
c_193 M10:DRN M8:GATE 8.30207e-19 
c_194 M10:DRN M9:DRN 2.8937e-20 
c_195 M10:DRN M9:GATE 4.58342e-18 
c_196 M10:DRN M9:SRC 1.97887e-17 
c_197 M10:DRN M10:GATE 3.43478e-17 
c_198 M10:DRN M11:DRN 8.34366e-19 
c_199 M10:DRN M11:GATE 1.44563e-18 
c_200 M10:DRN 0 8.36667e-18 
c_201 VDD M3:DRN 1.55542e-17 
c_202 VDD OE 8.15316e-17 
c_203 VDD M5:DRN 2.01732e-18 
c_204 VDD M1:DRN 3.53744e-17 
c_205 VDD M2:GATE 3.92768e-19 
c_206 VDD Z 3.78269e-17 
c_207 VDD M7:GATE 2.64016e-18 
c_208 VDD M8:GATE 1.02512e-17 
c_209 VDD M9:DRN 5.35094e-19 
c_210 VDD M9:GATE 1.01165e-17 
c_211 VDD M9:SRC 3.14133e-19 
c_212 VDD M10:GATE 7.53981e-18 
c_213 VDD M7:DRN 8.46473e-19 
c_214 VDD M11:DRN 2.91059e-17 
c_215 VDD M11:GATE 4.97107e-18 
c_216 VDD M12:SRC 2.07798e-18 
c_217 VDD M12:GATE 8.9745e-18 
c_218 VDD 0 1.15665e-16 
c_219 M12:DRN M1:GATE 2.02969e-17 
c_220 M12:DRN M2:GATE 5.70242e-19 
c_221 M12:DRN M2:SRC 1.0912e-20 
c_222 M12:DRN Z 8.13702e-19 
c_223 M12:DRN M9:DRN 1.14067e-21 
c_224 M12:DRN M9:SRC 1.1116e-19 
c_225 M12:DRN M10:GATE 2.79234e-18 
c_226 M12:DRN M11:DRN 1.82408e-17 
c_227 M12:DRN M11:GATE 2.58986e-17 
c_228 M12:DRN M12:SRC 6.71718e-19 
c_229 M12:DRN M12:GATE 2.66876e-17 
c_230 M12:DRN 0 1.30092e-17 
c_231 M8:DRN M3:DRN 2.96789e-18 
c_232 M8:DRN OE 3.93204e-18 
c_233 M8:DRN I:1 3.98983e-19 
c_234 M8:DRN M5:DRN 1.48291e-18 
c_235 M8:DRN M1:DRN 2.639e-20 
c_236 M8:DRN M2:SRC 5.40971e-20 
c_237 M8:DRN Z 2.19065e-19 
c_238 M8:DRN M7:GATE 2.71426e-17 
c_239 M8:DRN M8:GATE 3.10764e-17 
c_240 M8:DRN M9:DRN 6.52994e-18 
c_241 M8:DRN M9:GATE 1.02645e-17 
c_242 M8:DRN M9:SRC 9.10042e-18 
c_243 M8:DRN M10:GATE 5.58842e-18 
c_244 M8:DRN M7:DRN 1.83083e-18 
c_245 M8:DRN M11:DRN 1.0239e-17 
c_246 M8:DRN M11:GATE 4.36282e-18 
c_247 M8:DRN M12:SRC 9.19407e-18 
c_248 M8:DRN M12:GATE 4.3579e-18 
c_249 M8:DRN 0 7.25858e-17 

.ENDS
