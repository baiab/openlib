
.subckt CMPE32D1  A B CI S CO
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.06318p as=0.0567p l=0.09u nrd=0.298 nrs=0.268 pd=0.8955u ps=0.711u sa=3.726e-07 sb=1.161e-06 w=0.459u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.06723p as=0.06642p l=0.09u nrd=0.32 nrs=0.314 pd=0.918u ps=0.9081u sa=2.988e-07 sb=4.23e-07 w=0.459u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK nch ad=0.07128p as=0.05022p l=0.09u nrd=0.581 nrs=0.41 pd=1.17u ps=0.6939u sa=1.962e-07 sb=6.651e-07 w=0.351u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK nch ad=0.15714p as=0.06318p l=0.09u nrd=0.539 nrs=0.217 pd=1.926u ps=0.774u sa=1.3707e-06 sb=2.25e-07 w=0.54u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK nch ad=0.11178p as=0.0729p l=0.09u nrd=0.383 nrs=0.25 pd=1.494u ps=0.9675u sa=2.07e-07 sb=3.231e-07 w=0.54u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.07776p as=0.12636p l=0.09u nrd=0.266 nrs=0.433 pd=0.972u ps=1.548u sa=5.58e-07 sb=2.34e-07 w=0.54u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.11178p as=0.06399p l=0.09u nrd=0.383 nrs=0.22 pd=1.494u ps=0.936u sa=2.07e-07 sb=4.608e-07 w=0.54u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.06318p as=0.10368p l=0.09u nrd=0.217 nrs=0.357 pd=0.774u ps=1.782u sa=1.53e-07 sb=1.089e-06 w=0.54u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.06399p as=0.06318p l=0.09u nrd=0.22 nrs=0.217 pd=0.936u ps=0.774u sa=7.65e-07 sb=4.77e-07 w=0.54u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.03726p as=0.03969p l=0.09u nrd=0.507 nrs=0.543 pd=0.5265u ps=0.54u sa=9.036e-07 sb=1.503e-06 w=0.27u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK nch ad=0.06642p as=0.06399p l=0.09u nrd=0.227 nrs=0.22 pd=0.837u ps=0.936u sa=5.787e-07 sb=8.37e-07 w=0.54u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK nch ad=0.06399p as=0.06318p l=0.09u nrd=0.22 nrs=0.217 pd=0.936u ps=0.774u sa=9.819e-07 sb=5.49e-07 w=0.54u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK nch ad=0.04374p as=0.11178p l=0.09u nrd=0.417 nrs=1.065 pd=0.5805u ps=1.53u sa=5.31e-07 sb=2.25e-07 w=0.324u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.12636p as=0.07776p l=0.09u nrd=0.433 nrs=0.266 pd=1.548u ps=0.972u sa=2.34e-07 sb=5.58e-07 w=0.54u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.09477p as=0.06399p l=0.09u nrd=0.324 nrs=0.22 pd=1.512u ps=0.936u sa=4.95e-07 sb=1.701e-07 w=0.54u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.06318p as=0.06399p l=0.09u nrd=0.217 nrs=0.22 pd=0.774u ps=0.936u sa=4.77e-07 sb=7.65e-07 w=0.54u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.10368p as=0.06318p l=0.09u nrd=0.357 nrs=0.217 pd=1.782u ps=0.774u sa=1.089e-06 sb=1.53e-07 w=0.54u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK pch ad=0.12555p as=0.07209p l=0.09u nrd=0.341 nrs=0.196 pd=1.629u ps=0.873u sa=2.07e-07 sb=1.0179e-06 w=0.6075u 
MM30 M30:DRN M30:GATE M30:SRC M30:BULK pch ad=0.08424p as=0.08181p l=0.09u nrd=0.162 nrs=0.158 pd=0.954u ps=1.116u sa=4.77e-07 sb=7.65e-07 w=0.72u 
MM23 M23:DRN M23:GATE M23:SRC M23:BULK pch ad=0.14904p as=0.08586p l=0.09u nrd=0.287 nrs=0.166 pd=1.854u ps=1.125u sa=5.04e-07 sb=2.07e-07 w=0.72u 
MM32 M32:DRN M32:GATE M32:SRC M32:BULK pch ad=0.13122p as=0.08424p l=0.09u nrd=0.254 nrs=0.162 pd=2.142u ps=0.954u sa=1.089e-06 sb=1.53e-07 w=0.72u 
MM25 M25:DRN M25:GATE M25:SRC M25:BULK pch ad=0.09072p as=0.11907p l=0.09u nrd=0.175 nrs=0.23 pd=0.972u ps=1.197u sa=9.414e-07 sb=8.46e-07 w=0.72u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK pch ad=0.11016p as=0.0648p l=0.09u nrd=0.39 nrs=0.23 pd=1.476u ps=0.8343u sa=4.608e-07 sb=2.07e-07 w=0.531u 
MM34 M34:DRN M34:GATE M34:SRC M34:BULK pch ad=0.14904p as=0.08586p l=0.09u nrd=0.287 nrs=0.166 pd=1.854u ps=1.125u sa=2.07e-07 sb=5.04e-07 w=0.72u 
MM27 M27:DRN M27:GATE M27:SRC M27:BULK pch ad=0.11907p as=0.08424p l=0.09u nrd=0.23 nrs=0.162 pd=1.197u ps=0.954u sa=1.3824e-06 sb=4.77e-07 w=0.72u 
MM29 M29:DRN M29:GATE M29:SRC M29:BULK pch ad=0.09882p as=0.16848p l=0.09u nrd=0.19 nrs=0.325 pd=1.152u ps=1.908u sa=5.274e-07 sb=2.34e-07 w=0.72u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK pch ad=0.14175p as=0.08343p l=0.09u nrd=0.303 nrs=0.178 pd=1.782u ps=1.0737u sa=2.07e-07 sb=3.231e-07 w=0.684u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK pch ad=0.08586p as=0.08748p l=0.09u nrd=0.166 nrs=0.168 pd=1.035u ps=1.1061u sa=3.915e-07 sb=4.986e-07 w=0.72u 
MM31 M31:DRN M31:GATE M31:SRC M31:BULK pch ad=0.08424p as=0.13122p l=0.09u nrd=0.162 nrs=0.254 pd=0.954u ps=2.142u sa=1.53e-07 sb=1.089e-06 w=0.72u 
MM24 M24:DRN M24:GATE M24:SRC M24:BULK pch ad=0.08748p as=0.09072p l=0.09u nrd=0.168 nrs=0.175 pd=1.1061u ps=0.972u sa=4.302e-07 sb=1.188e-06 w=0.72u 
MM33 M33:DRN M33:GATE M33:SRC M33:BULK pch ad=0.08181p as=0.08424p l=0.09u nrd=0.158 nrs=0.162 pd=1.116u ps=0.954u sa=7.65e-07 sb=4.77e-07 w=0.72u 
MM26 M26:DRN M26:GATE M26:SRC M26:BULK pch ad=0.14823p as=0.08424p l=0.09u nrd=0.287 nrs=0.162 pd=2.322u ps=0.954u sa=1.7406e-06 sb=1.53e-07 w=0.72u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK pch ad=0.06318p as=0.06318p l=0.09u nrd=0.232 nrs=0.232 pd=0.8019u ps=0.8019u sa=7.29e-07 sb=1.512e-06 w=0.522u 
MM28 M28:DRN M28:GATE M28:SRC M28:BULK pch ad=0.14742p as=0.09882p l=0.09u nrd=0.285 nrs=0.19 pd=1.908u ps=1.152u sa=2.007e-07 sb=5.58e-07 w=0.72u 
R1 M20:DRN M8:SRC 57.3338
R2 M20:DRN M16:DRN 55.086
R3 M20:DRN M32:SRC 101.28
R4 M32:SRC M8:SRC 58.5711
R5 M32:SRC M16:DRN 56.2749
R6 M32:SRC M33:SRC 0.001
R7 M8:SRC M16:DRN 27.3389
R8 M8:SRC M7:SRC 0.001
R9 M4:SRC M3:SRC 0.001
R10 M4:SRC M7:DRN 1.36364e-09
R11 M17:BULK M6:SRC 7.93854e-06
R12 M17:BULK M7:DRN 0.000857339
R13 M17:BULK M16:BULK 0.001
R14 M17:BULK M4:BULK 0.001
R15 M17:BULK M6:BULK 0.001
R16 M17:BULK M5:BULK 0.001
R17 M17:BULK M8:BULK 0.001
R18 M17:BULK M7:BULK 0.001
R19 M17:BULK M3:BULK 0.001
R20 M17:BULK M12:BULK 0.001
R21 M17:BULK M10:BULK 0.001
R22 M17:BULK M11:BULK 0.001
R23 M17:BULK M9:BULK 0.001
R24 M17:BULK M13:BULK 0.001
R25 M17:BULK M15:BULK 0.001
R26 M17:BULK M14:BULK 0.001
R27 M17:BULK M1:BULK 0.001
R28 M17:BULK M2:BULK 0.001
R29 GND:1 M6:SRC 49.6834
R30 GND:1 M7:DRN 1.15959
R31 GND:1 GND 1.17912
R32 GND:1 M14:DRN 18
R33 GND:1 M2:DRN 19.2357
R34 GND M6:SRC 4.14797
R35 GND M7:DRN 2.9389
R36 M14:DRN M7:DRN 8e-10
R37 M13:SRC M7:DRN 1.83333e-09
R38 M13:SRC M15:DRN 0.001
R39 M2:DRN M7:DRN 1.11538e-09
R40 M2:DRN M1:SRC 0.001
R41 M6:SRC M7:DRN 1.36517e-09
R42 M6:SRC M5:SRC 9.90741e-10
R43 M5:SRC M8:DRN 0.001
R44 M29:SRC S 9.29909
R45 S M2:SRC 9.20846
R46 M28:DRN CO 18.2296
R47 CO M1:DRN 9.22277
R48 M25:DRN M13:DRN 36.5011
R49 M25:DRN M24:SRC 0.001
R50 M13:DRN M9:SRC 1.0641e-09
R51 M29:GATE N_20:1 91.162
R52 M29:GATE M2:GATE 275.474
R53 M24:DRN N_20:1 18
R54 M24:DRN M19:SRC 0.001
R55 N_20:1 M11:DRN 18.685
R56 N_20:1 M2:GATE 87.6003
R57 M11:DRN M9:DRN 0.001
R58 M28:GATE M22:DRN 209.779
R59 M28:GATE M12:SRC 437.678
R60 M28:GATE M1:GATE 123.12
R61 M22:DRN M12:SRC 28.8773
R62 M22:DRN M21:SRC 0.001
R63 M12:SRC M10:SRC 0.001
R64 M24:GATE M11:GATE 134.4
R65 M24:GATE M22:GATE 186.84
R66 M22:GATE M3:DRN 554.475
R67 M22:GATE M12:GATE 188.581
R68 M22:GATE M23:DRN 555.4
R69 M23:DRN M3:DRN 40.5039
R70 M23:DRN M12:GATE 280.209
R71 M12:GATE M3:DRN 279.742
R72 M34:GATE M4:GATE 313.965
R73 M34:GATE B 88.7579
R74 M34:GATE M20:GATE 223.56
R75 B M4:GATE 82.0872
R76 M4:GATE M17:GATE 154.92
R77 N_17:1 M8:GATE 48.16
R78 N_17:1 N_17:3 16.2972
R79 N_17:1 M33:GATE 65.88
R80 N_17:1 N_17:2 12.5545
R81 N_17:1 M6:DRN 770.973
R82 N_17:2 M7:GATE 48.16
R83 N_17:2 N_17:3 16.4613
R84 N_17:2 M32:GATE 65.88
R85 N_17:2 M6:DRN 778.735
R86 N_17:3 M17:SRC 25.3258
R87 N_17:3 M18:DRN 12.0281
R88 N_17:3 M31:DRN 9.1017
R89 N_17:3 M6:DRN 9.65402
R90 M31:DRN M18:DRN 1177.4
R91 M31:DRN M30:DRN 0.001
R92 M18:DRN M17:SRC 110.984
R93 M6:DRN M5:DRN 0.001
R94 N_24:1 M16:SRC 301.904
R95 N_24:1 M20:SRC 317.753
R96 N_24:1 M3:GATE 270.143
R97 N_24:1 M9:GATE 130.2
R98 N_24:1 M10:GATE 42.72
R99 M21:GATE M23:GATE 177.84
R100 M23:GATE M3:GATE 121.942
R101 M19:GATE M10:GATE 133.309
R102 M3:GATE M16:SRC 290.961
R103 M3:GATE M20:SRC 306.236
R104 M20:SRC M16:SRC 42.0539
R105 M20:SRC M18:SRC 0.001
R106 M17:DRN M16:SRC 0.001
R107 A:1 M30:GATE 105.704
R108 A:1 A 21.8465
R109 A:1 M5:GATE 88.655
R110 A:1 M6:GATE 56.16
R111 A:1 M31:GATE 66.96
R112 M30:GATE M5:GATE 335.904
R113 N_12:1 M16:GATE 117.615
R114 N_12:1 M34:DRN 9.18055
R115 N_12:1 M4:DRN 18.6916
R116 N_12:1 M12:DRN 22.2095
R117 N_12:1 M18:GATE 87.548
R118 N_12:1 M21:DRN 10.6216
R119 M34:DRN M21:DRN 633.156
R120 M21:DRN M12:DRN 188.382
R121 M4:DRN M16:GATE 6966.39
R122 M4:DRN M18:GATE 5185.51
R123 M18:GATE M16:GATE 448.945
R124 CI:1 M15:GATE 43.84
R125 CI:1 CI 10.4629
R126 CI:1 M14:GATE 99.096
R127 CI:1 M27:GATE 70.2
R128 CI:1 M26:GATE 160.821
R129 M26:GATE CI 194.865
R130 M26:GATE M14:GATE 558.24
R131 CI M14:GATE 120.074
R132 N_5:1 M13:GATE 67.9904
R133 N_5:1 M11:SRC 24.4794
R134 N_5:1 M27:SRC 18
R135 N_5:1 M14:SRC 21.5731
R136 N_5:1 M22:SRC 25.2138
R137 N_5:1 M25:GATE 106.211
R138 M25:GATE M13:GATE 290.081
R139 M22:SRC M11:SRC 172.885
R140 M22:SRC M14:SRC 347.635
R141 M22:SRC M19:DRN 0.001
R142 M27:SRC M26:SRC 0.001
R143 M14:SRC M11:SRC 337.509
R144 M14:SRC M15:SRC 0.001
R145 M11:SRC M10:DRN 0.001
R146 VDD:1 M31:SRC 20.7127
R147 VDD:1 VDD 0.499816
R148 VDD:1 M34:SRC 2.42887
R149 VDD:1 M32:DRN 4.40523
R150 VDD:1 VDD:2 0.687437
R151 VDD:2 M34:SRC 2.01006
R152 VDD:2 M25:SRC 19.533
R153 VDD:2 M28:SRC 18.1179
R154 M34:BULK M31:SRC 7.8626e-06
R155 M34:BULK M34:SRC 0.00474834
R156 M34:BULK M30:SRC 0.00514403
R157 M34:BULK M32:DRN 0.00514403
R158 M34:BULK M23:BULK 0.001
R159 M34:BULK M25:SRC 0.00293945
R160 M34:BULK M26:DRN 0.00280584
R161 M34:BULK M28:SRC 0.00385802
R162 M34:BULK M21:BULK 0.001
R163 M34:BULK M31:BULK 0.001
R164 M34:BULK M30:BULK 0.001
R165 M34:BULK M33:BULK 0.001
R166 M34:BULK M32:BULK 0.001
R167 M34:BULK M20:BULK 0.001
R168 M34:BULK M18:BULK 0.001
R169 M34:BULK M22:BULK 0.001
R170 M34:BULK M19:BULK 0.001
R171 M34:BULK M24:BULK 0.001
R172 M34:BULK M25:BULK 0.001
R173 M34:BULK M27:BULK 0.001
R174 M34:BULK M26:BULK 0.001
R175 M34:BULK M28:BULK 0.001
R176 M34:BULK M29:BULK 0.001
R177 M34:SRC M32:DRN 1.42222e-09
R178 M34:SRC M25:SRC 5.71429e-10
R179 M34:SRC M26:DRN 0.001
R180 M34:SRC M28:SRC 4.60714e-10
R181 M34:SRC M23:SRC 0.001
R182 M25:SRC M27:DRN 0.001
R183 M28:SRC M29:DRN 0.001
R184 VDD M31:SRC 4.46006
R185 VDD M32:DRN 10.3408
R186 M31:SRC M30:SRC 1e-09
R187 M31:SRC M32:DRN 1.35e-09
R188 M30:SRC M33:DRN 0.001
c_1 M20:DRN 0 5.60421e-18 
c_2 M32:SRC 0 2.41597e-17 
c_3 M8:SRC 0 2.73394e-19 
c_4 M16:DRN 0 4.20856e-18 
c_5 M4:SRC 0 3.2646e-18 
c_6 M17:BULK M8:SRC 1.01413e-17 
c_7 M17:BULK 0 2.71383e-17 
c_8 GND:1 M8:SRC 2.12457e-18 
c_9 GND:1 M16:DRN 2.11197e-17 
c_10 GND:1 M32:SRC 7.25709e-17 
c_11 GND:1 0 2.44816e-16 
c_12 GND 0 7.34585e-18 
c_13 M14:DRN 0 2.28279e-18 
c_14 M13:SRC 0 3.03795e-18 
c_15 M2:DRN 0 6.16044e-18 
c_16 M6:SRC M8:SRC 1.11888e-17 
c_17 M6:SRC M16:DRN 1.00533e-17 
c_18 M6:SRC M32:SRC 4.42193e-20 
c_19 M6:SRC 0 2.05122e-16 
c_20 M5:SRC M16:DRN 6.85193e-20 
c_21 M5:SRC 0 4.1912e-18 
c_22 M7:DRN M16:DRN 3.54719e-17 
c_23 M7:DRN 0 3.80816e-17 
c_24 M29:SRC M6:SRC 3.55798e-20 
c_25 M29:SRC 0 6.59337e-18 
c_26 S M6:SRC 9.64926e-20 
c_27 S M7:DRN 1.16423e-18 
c_28 S M17:BULK 2.94231e-18 
c_29 S GND:1 7.82837e-17 
c_30 S M2:DRN 2.52378e-19 
c_31 S 0 5.31825e-17 
c_32 M2:SRC M6:SRC 1.02089e-17 
c_33 M2:SRC M7:DRN 1.5674e-18 
c_34 M2:SRC GND:1 1.87328e-18 
c_35 M2:SRC M2:DRN 9.81276e-19 
c_36 M2:SRC 0 2.70517e-18 
c_37 M28:DRN M6:SRC 3.55798e-20 
c_38 M28:DRN 0 3.47329e-18 
c_39 CO M6:SRC 1.38364e-19 
c_40 CO M7:DRN 1.76778e-18 
c_41 CO M17:BULK 2.03352e-18 
c_42 CO GND:1 8.47685e-17 
c_43 CO M14:DRN 1.81694e-20 
c_44 CO M2:DRN 6.03506e-19 
c_45 CO 0 2.23527e-17 
c_46 M1:DRN M6:SRC 1.02089e-17 
c_47 M1:DRN M7:DRN 1.68451e-18 
c_48 M1:DRN GND:1 2.91778e-18 
c_49 M1:DRN M14:DRN 2.94867e-17 
c_50 M1:DRN M2:DRN 5.71396e-19 
c_51 M1:DRN 0 5.13857e-18 
c_52 M25:DRN M6:SRC 8.21131e-20 
c_53 M25:DRN M7:DRN 6.64033e-19 
c_54 M25:DRN M17:BULK 2.12037e-18 
c_55 M25:DRN 0 1.99327e-17 
c_56 M13:DRN M6:SRC 1.12438e-18 
c_57 M13:DRN M7:DRN 2.34433e-19 
c_58 M13:DRN GND:1 1.60956e-18 
c_59 M13:DRN 0 1.3037e-17 
c_60 M9:SRC M6:SRC 8.26669e-18 
c_61 M29:GATE M2:SRC 1.05082e-17 
c_62 M29:GATE S 1.78469e-17 
c_63 M29:GATE M28:DRN 1.06341e-19 
c_64 M29:GATE M29:SRC 3.55592e-17 
c_65 M29:GATE 0 9.04628e-18 
c_66 M24:DRN M6:SRC 7.81031e-20 
c_67 M24:DRN M7:DRN 7.51825e-24 
c_68 M24:DRN M25:DRN 1.77119e-19 
c_69 M24:DRN CO 1.04638e-19 
c_70 N_20:1 M6:SRC 3.81138e-21 
c_71 N_20:1 M7:DRN 1.68889e-17 
c_72 N_20:1 M17:BULK 7.84415e-18 
c_73 N_20:1 GND:1 2.69262e-17 
c_74 N_20:1 M25:DRN 7.34472e-17 
c_75 N_20:1 M13:DRN 4.057e-17 
c_76 N_20:1 M14:DRN 1.35343e-19 
c_77 N_20:1 CO 7.60426e-17 
c_78 N_20:1 M1:DRN 4.1146e-20 
c_79 N_20:1 M2:DRN 1.51916e-18 
c_80 N_20:1 M2:SRC 1.26086e-19 
c_81 N_20:1 S 9.60713e-17 
c_82 N_20:1 M28:DRN 6.6792e-18 
c_83 N_20:1 M29:SRC 1.16621e-18 
c_84 N_20:1 0 1.9726e-17 
c_85 M2:GATE M6:SRC 4.3585e-18 
c_86 M2:GATE M7:DRN 1.69718e-17 
c_87 M2:GATE M17:BULK 1.20737e-18 
c_88 M2:GATE GND:1 6.92465e-18 
c_89 M2:GATE M14:DRN 1.19929e-19 
c_90 M2:GATE M2:DRN 2.16574e-17 
c_91 M2:GATE M2:SRC 2.47358e-17 
c_92 M2:GATE S 1.20935e-17 
c_93 M11:DRN M6:SRC 6.5597e-18 
c_94 M11:DRN M7:DRN 2.0292e-20 
c_95 M11:DRN GND:1 3.17901e-18 
c_96 M11:DRN M25:DRN 1.2256e-18 
c_97 M11:DRN M13:DRN 1.06905e-18 
c_98 M11:DRN M13:SRC 7.77571e-20 
c_99 M11:DRN M28:DRN 4.12496e-19 
c_100 M11:DRN 0 4.7931e-19 
c_101 M28:GATE M6:SRC 2.95674e-19 
c_102 M28:GATE M7:DRN 9.66998e-19 
c_103 M28:GATE M17:BULK 3.85165e-18 
c_104 M28:GATE GND:1 6.70861e-18 
c_105 M28:GATE N_20:1 1.90066e-17 
c_106 M28:GATE M11:DRN 1.30623e-19 
c_107 M28:GATE CO 1.00121e-17 
c_108 M28:GATE M1:DRN 7.57706e-18 
c_109 M28:GATE M2:DRN 1.21461e-17 
c_110 M28:GATE M29:GATE 7.01269e-18 
c_111 M28:GATE 0 1.82577e-17 
c_112 M22:DRN M6:SRC 3.58804e-20 
c_113 M22:DRN M7:DRN 1.3318e-19 
c_114 M22:DRN M17:BULK 4.6002e-18 
c_115 M22:DRN N_20:1 2.20213e-16 
c_116 M22:DRN M24:DRN 3.15242e-18 
c_117 M22:DRN M14:DRN 1.10115e-18 
c_118 M22:DRN 0 3.11957e-19 
c_119 M1:GATE M6:SRC 4.3585e-18 
c_120 M1:GATE M7:DRN 3.56782e-17 
c_121 M1:GATE M17:BULK 4.03786e-18 
c_122 M1:GATE GND:1 3.86811e-18 
c_123 M1:GATE N_20:1 2.04297e-17 
c_124 M1:GATE M14:DRN 1.38369e-18 
c_125 M1:GATE CO 5.10942e-18 
c_126 M1:GATE M1:DRN 2.59603e-17 
c_127 M1:GATE M2:DRN 6.36218e-18 
c_128 M1:GATE M2:GATE 2.37049e-18 
c_129 M1:GATE 0 4.10197e-19 
c_130 M12:SRC M6:SRC 7.54651e-18 
c_131 M12:SRC M7:DRN 3.45713e-20 
c_132 M12:SRC GND:1 2.28655e-17 
c_133 M12:SRC M4:SRC 2.88336e-21 
c_134 M12:SRC M11:DRN 1.13047e-19 
c_135 M12:SRC M13:SRC 1.66989e-22 
c_136 M12:SRC CO 5.88458e-18 
c_137 M12:SRC M28:DRN 4.27227e-17 
c_138 M12:SRC M29:GATE 2.35393e-18 
c_139 M12:SRC 0 2.9817e-17 
c_140 M24:GATE M22:DRN 2.0347e-17 
c_141 M24:GATE M12:SRC 3.89111e-19 
c_142 M24:GATE N_20:1 8.63544e-18 
c_143 M24:GATE M11:DRN 1.43097e-20 
c_144 M24:GATE 0 6.78016e-18 
c_145 M22:GATE M22:DRN 6.23756e-17 
c_146 M22:GATE M24:DRN 1.49719e-17 
c_147 M22:GATE 0 1.49772e-17 
c_148 M23:DRN M22:DRN 4.60704e-19 
c_149 M23:DRN 0 3.80433e-18 
c_150 M12:GATE M22:DRN 4.49271e-18 
c_151 M12:GATE M12:SRC 3.1884e-17 
c_152 M12:GATE 0 1.9372e-17 
c_153 M11:GATE M22:DRN 4.61338e-20 
c_154 M11:GATE M25:DRN 1.91361e-17 
c_155 M11:GATE N_20:1 1.84584e-17 
c_156 M11:GATE M11:DRN 3.3042e-17 
c_157 M11:GATE M24:DRN 2.76164e-17 
c_158 M11:GATE M13:DRN 3.35344e-18 
c_159 M11:GATE 0 2.10605e-18 
c_160 M3:DRN M22:DRN 1.78322e-20 
c_161 M3:DRN M12:SRC 2.54749e-19 
c_162 M3:DRN 0 1.09757e-17 
c_163 M34:GATE M3:DRN 4.96269e-19 
c_164 M34:GATE M4:SRC 2.60665e-18 
c_165 M34:GATE M20:DRN 2.90382e-18 
c_166 M34:GATE M23:DRN 1.274e-19 
c_167 M34:GATE 0 4.32052e-18 
c_168 B M6:SRC 5.71707e-20 
c_169 B M7:DRN 7.94503e-19 
c_170 B M17:BULK 6.68816e-18 
c_171 B M3:DRN 6.63692e-17 
c_172 B M12:GATE 2.30914e-19 
c_173 B GND:1 2.51833e-19 
c_174 B M4:SRC 1.23172e-18 
c_175 B M23:DRN 1.52891e-19 
c_176 B 0 2.47578e-19 
c_177 M4:GATE M7:DRN 7.06972e-18 
c_178 M4:GATE M17:BULK 2.27587e-18 
c_179 M4:GATE M3:DRN 1.11439e-18 
c_180 M4:GATE M12:GATE 1.008e-19 
c_181 M4:GATE GND:1 1.13153e-18 
c_182 M4:GATE 0 2.80415e-19 
c_183 M20:GATE M8:SRC 6.79717e-18 
c_184 M20:GATE M20:DRN 1.67703e-17 
c_185 M20:GATE M24:GATE 1.60224e-20 
c_186 M20:GATE M32:SRC 1.11479e-20 
c_187 M20:GATE 0 8.86156e-19 
c_188 M17:GATE M6:SRC 3.03456e-17 
c_189 M17:GATE M8:SRC 4.92585e-19 
c_190 M17:GATE M7:DRN 4.22145e-17 
c_191 M17:GATE M16:DRN 8.25538e-20 
c_192 M17:GATE M17:BULK 7.8284e-18 
c_193 M17:GATE M3:DRN 9.97742e-19 
c_194 M17:GATE M12:GATE 2.4669e-21 
c_195 M17:GATE GND:1 2.59755e-17 
c_196 M17:GATE 0 1.6146e-20 
c_197 N_17:1 M6:SRC 7.02512e-20 
c_198 N_17:1 M8:SRC 3.97427e-17 
c_199 N_17:1 M16:DRN 8.61435e-18 
c_200 N_17:1 M17:BULK 5.27718e-18 
c_201 N_17:1 GND:1 6.36112e-19 
c_202 N_17:1 B 3.29317e-21 
c_203 N_17:1 M32:SRC 1.52529e-17 
c_204 N_17:1 M20:GATE 4.34712e-19 
c_205 N_17:1 0 5.83062e-18 
c_206 N_17:2 M8:SRC 3.26121e-17 
c_207 N_17:2 M16:DRN 2.26109e-18 
c_208 N_17:2 M17:BULK 2.94701e-18 
c_209 N_17:2 GND:1 5.73667e-19 
c_210 N_17:2 B 2.08847e-20 
c_211 N_17:2 M20:GATE 7.59746e-19 
c_212 N_17:2 0 5.95362e-18 
c_213 N_17:3 M6:SRC 1.50129e-18 
c_214 N_17:3 M8:SRC 2.30798e-17 
c_215 N_17:3 M7:DRN 1.18706e-18 
c_216 N_17:3 M16:DRN 1.2067e-16 
c_217 N_17:3 M17:BULK 9.95088e-18 
c_218 N_17:3 GND:1 4.82349e-17 
c_219 N_17:3 M20:DRN 8.81973e-17 
c_220 N_17:3 M5:SRC 4.04257e-18 
c_221 N_17:3 M32:SRC 6.83264e-18 
c_222 N_17:3 M20:GATE 1.12844e-17 
c_223 N_17:3 0 1.25234e-18 
c_224 M33:GATE M16:DRN 5.48644e-18 
c_225 M33:GATE M34:GATE 2.45016e-20 
c_226 M33:GATE M20:DRN 1.11479e-20 
c_227 M33:GATE M32:SRC 1.69133e-17 
c_228 M33:GATE M20:GATE 4.61739e-20 
c_229 M33:GATE 0 2.51152e-20 
c_230 M32:GATE M8:SRC 1.09994e-17 
c_231 M32:GATE M34:GATE 2.3362e-19 
c_232 M32:GATE B 2.25548e-23 
c_233 M32:GATE M20:DRN 1.83381e-18 
c_234 M32:GATE M32:SRC 1.67633e-17 
c_235 M32:GATE M20:GATE 1.16869e-18 
c_236 M32:GATE 0 2.1803e-18 
c_237 M31:DRN M6:SRC 4.42193e-20 
c_238 M31:DRN M16:DRN 3.47664e-20 
c_239 M31:DRN M32:SRC 5.78741e-20 
c_240 M31:DRN 0 4.35054e-18 
c_241 M18:DRN M17:GATE 4.66334e-18 
c_242 M18:DRN M6:SRC 4.49724e-21 
c_243 M18:DRN B 8.23008e-19 
c_244 M18:DRN M20:DRN 7.14018e-19 
c_245 M18:DRN M20:GATE 6.75275e-18 
c_246 M7:GATE M17:GATE 2.17955e-19 
c_247 M7:GATE M6:SRC 9.11383e-18 
c_248 M7:GATE M8:SRC 1.27657e-18 
c_249 M7:GATE M7:DRN 1.39247e-17 
c_250 M7:GATE M16:DRN 1.4326e-17 
c_251 M7:GATE M17:BULK 3.13373e-18 
c_252 M7:GATE GND:1 4.93541e-18 
c_253 M7:GATE M5:SRC 9.89998e-19 
c_254 M7:GATE 0 6.58889e-19 
c_255 M8:GATE M17:GATE 1.98564e-21 
c_256 M8:GATE M6:SRC 9.4454e-18 
c_257 M8:GATE M8:SRC 1.13044e-17 
c_258 M8:GATE M7:DRN 1.51356e-18 
c_259 M8:GATE M16:DRN 4.60206e-18 
c_260 M8:GATE M17:BULK 4.6675e-18 
c_261 M8:GATE GND:1 1.03078e-18 
c_262 M8:GATE M5:SRC 1.03026e-17 
c_263 M8:GATE 0 1.18309e-18 
c_264 M6:DRN M6:SRC 1.1194e-17 
c_265 M6:DRN M8:SRC 4.34055e-20 
c_266 M6:DRN GND:1 2.22919e-18 
c_267 M6:DRN 0 5.57119e-18 
c_268 M17:SRC M17:GATE 1.58775e-17 
c_269 M17:SRC M6:SRC 6.99815e-18 
c_270 M17:SRC M8:SRC 5.91914e-19 
c_271 M17:SRC M7:DRN 3.58216e-20 
c_272 M17:SRC M16:DRN 9.61698e-19 
c_273 M17:SRC M4:GATE 1.78363e-17 
c_274 M17:SRC GND:1 2.87418e-18 
c_275 M17:SRC M34:GATE 4.22355e-18 
c_276 M17:SRC M4:SRC 4.34055e-20 
c_277 M17:SRC B 1.07993e-18 
c_278 M17:SRC 0 1.637e-17 
c_279 N_24:1 M7:DRN 6.21854e-20 
c_280 N_24:1 M17:BULK 4.13081e-18 
c_281 N_24:1 M12:GATE 2.45947e-18 
c_282 N_24:1 GND:1 1.00281e-16 
c_283 N_24:1 M22:DRN 4.37125e-18 
c_284 N_24:1 M12:SRC 1.59791e-17 
c_285 N_24:1 M11:GATE 6.49258e-19 
c_286 N_24:1 M11:DRN 1.34722e-17 
c_287 N_24:1 M13:DRN 8.35079e-18 
c_288 N_24:1 M13:SRC 9.64391e-19 
c_289 N_24:1 0 9.4184e-18 
c_290 M21:GATE M4:GATE 1.5844e-20 
c_291 M21:GATE M3:DRN 8.03706e-19 
c_292 M21:GATE M12:GATE 5.59956e-18 
c_293 M21:GATE N_17:3 2.24828e-19 
c_294 M21:GATE M34:GATE 3.58271e-20 
c_295 M21:GATE M22:DRN 2.56331e-17 
c_296 M21:GATE M23:DRN 1.71346e-17 
c_297 M21:GATE M24:GATE 1.85197e-19 
c_298 M21:GATE M20:GATE 1.30674e-20 
c_299 M21:GATE M22:GATE 5.05565e-18 
c_300 M23:GATE M6:SRC 2.27042e-20 
c_301 M23:GATE M7:DRN 7.84274e-21 
c_302 M23:GATE M17:BULK 4.36238e-18 
c_303 M23:GATE M17:SRC 1.6948e-19 
c_304 M23:GATE M18:DRN 6.49973e-21 
c_305 M23:GATE M3:DRN 1.07019e-21 
c_306 M23:GATE M12:GATE 1.45597e-19 
c_307 M23:GATE M34:GATE 2.47912e-17 
c_308 M23:GATE M4:SRC 5.02015e-19 
c_309 M23:GATE B 1.02807e-17 
c_310 M23:GATE M22:DRN 1.81798e-17 
c_311 M23:GATE M32:GATE 2.82272e-21 
c_312 M23:GATE M23:DRN 6.02162e-18 
c_313 M23:GATE M24:GATE 3.0584e-18 
c_314 M23:GATE M20:GATE 1.49191e-18 
c_315 M23:GATE M22:GATE 2.47465e-18 
c_316 M19:GATE M7:DRN 1.96357e-21 
c_317 M19:GATE M17:BULK 5.10014e-18 
c_318 M19:GATE M12:GATE 5.21955e-18 
c_319 M19:GATE GND:1 4.3718e-20 
c_320 M19:GATE N_17:3 8.67649e-20 
c_321 M19:GATE M22:DRN 1.01254e-17 
c_322 M19:GATE M12:SRC 4.78526e-18 
c_323 M19:GATE M24:GATE 6.62025e-18 
c_324 M19:GATE M25:DRN 6.58791e-20 
c_325 M19:GATE N_20:1 1.33796e-19 
c_326 M19:GATE M11:DRN 2.24334e-19 
c_327 M19:GATE M24:DRN 5.88026e-18 
c_328 M19:GATE M22:GATE 1.75018e-17 
c_329 M19:GATE 0 2.21594e-18 
c_330 M3:GATE M6:SRC 7.03594e-17 
c_331 M3:GATE M7:GATE 6.27271e-22 
c_332 M3:GATE M7:DRN 4.5311e-17 
c_333 M3:GATE M17:BULK 8.95288e-18 
c_334 M3:GATE M17:SRC 4.23265e-20 
c_335 M3:GATE M4:GATE 8.69267e-18 
c_336 M3:GATE M12:GATE 1.60458e-17 
c_337 M3:GATE GND:1 5.64701e-17 
c_338 M3:GATE M23:DRN 3.94318e-17 
c_339 M3:GATE M12:SRC 1.61665e-17 
c_340 M3:GATE M11:GATE 4.63962e-18 
c_341 M3:GATE M13:SRC 1.08638e-18 
c_342 M3:GATE M22:GATE 1.12552e-20 
c_343 M3:GATE 0 1.33909e-19 
c_344 M9:GATE M7:DRN 5.26184e-20 
c_345 M9:GATE M17:BULK 6.01142e-18 
c_346 M9:GATE M25:DRN 8.00321e-18 
c_347 M9:GATE M11:GATE 1.03971e-17 
c_348 M9:GATE N_20:1 4.22387e-18 
c_349 M9:GATE M11:DRN 1.87828e-17 
c_350 M9:GATE M13:DRN 1.16758e-17 
c_351 M9:GATE M9:SRC 1.96123e-18 
c_352 M9:GATE 0 2.59937e-18 
c_353 M10:GATE GND:1 6.26987e-19 
c_354 M10:GATE M24:GATE 2.29268e-17 
c_355 M10:GATE M24:DRN 1.66446e-17 
c_356 M10:GATE N_20:1 8.2391e-18 
c_357 M10:GATE M11:GATE 3.93761e-18 
c_358 M10:GATE 0 5.40454e-18 
c_359 M20:SRC M17:GATE 2.7734e-17 
c_360 M20:SRC M6:SRC 4.49724e-21 
c_361 M20:SRC M8:SRC 6.41102e-18 
c_362 M20:SRC M17:BULK 1.18082e-17 
c_363 M20:SRC M17:SRC 4.34421e-18 
c_364 M20:SRC M18:DRN 1.20415e-18 
c_365 M20:SRC M4:GATE 6.55001e-18 
c_366 M20:SRC M3:DRN 9.61386e-17 
c_367 M20:SRC M12:GATE 3.29433e-18 
c_368 M20:SRC GND:1 7.94656e-17 
c_369 M20:SRC N_17:3 4.39489e-18 
c_370 M20:SRC M34:GATE 1.49415e-17 
c_371 M20:SRC M4:SRC 4.18463e-18 
c_372 M20:SRC B 7.86849e-18 
c_373 M20:SRC M22:DRN 5.76614e-18 
c_374 M20:SRC M32:GATE 1.11479e-20 
c_375 M20:SRC M20:DRN 4.28173e-19 
c_376 M20:SRC M32:SRC 9.99407e-22 
c_377 M20:SRC M20:GATE 2.70296e-17 
c_378 M20:SRC N_20:1 9.69636e-19 
c_379 M20:SRC M24:DRN 1.8231e-19 
c_380 M20:SRC M14:DRN 7.46845e-21 
c_381 M20:SRC 0 2.17045e-19 
c_382 M17:DRN M7:DRN 3.94267e-20 
c_383 M17:DRN M6:SRC 8.11352e-18 
c_384 M17:DRN M17:SRC 7.9311e-18 
c_385 M17:DRN M17:GATE 1.025e-17 
c_386 M16:SRC M17:GATE 1.89594e-17 
c_387 M16:SRC M6:SRC 2.37052e-18 
c_388 M16:SRC M8:SRC 1.19118e-16 
c_389 M16:SRC M7:GATE 1.03701e-20 
c_390 M16:SRC M7:DRN 7.2637e-17 
c_391 M16:SRC M16:DRN 2.62881e-18 
c_392 M16:SRC M18:DRN 3.18482e-19 
c_393 M16:SRC M4:GATE 1.62172e-19 
c_394 M16:SRC GND:1 2.55549e-18 
c_395 M16:SRC N_17:3 1.76662e-16 
c_396 M16:SRC M31:DRN 1.60073e-19 
c_397 M16:SRC N_17:1 5.69368e-19 
c_398 M16:SRC M33:GATE 1.96047e-19 
c_399 M16:SRC N_17:2 2.08859e-19 
c_400 M16:SRC M32:GATE 2.84126e-19 
c_401 M16:SRC M20:DRN 1.72153e-18 
c_402 M16:SRC M23:DRN 8.68086e-21 
c_403 M16:SRC M12:SRC 6.44718e-21 
c_404 M16:SRC M24:GATE 1.35577e-19 
c_405 M16:SRC M25:DRN 5.93473e-21 
c_406 M16:SRC 0 1.82252e-19 
c_407 A:1 M6:SRC 8.41684e-18 
c_408 A:1 M17:BULK 8.32718e-18 
c_409 A:1 GND:1 1.19115e-18 
c_410 A:1 N_17:3 1.02542e-17 
c_411 A:1 M31:DRN 7.5221e-18 
c_412 A:1 N_17:1 3.43352e-19 
c_413 A:1 M6:DRN 7.90492e-17 
c_414 A:1 GND 7.22942e-21 
c_415 A:1 0 4.01428e-20 
c_416 M31:GATE N_17:3 1.23595e-17 
c_417 M31:GATE M33:GATE 3.71892e-19 
c_418 M31:GATE M31:DRN 3.37538e-17 
c_419 M31:GATE 0 5.55772e-19 
c_420 M30:GATE M17:BULK 2.93209e-18 
c_421 M30:GATE N_17:3 1.18549e-17 
c_422 M30:GATE M31:DRN 3.38357e-17 
c_423 M30:GATE N_17:1 2.58198e-18 
c_424 M30:GATE M33:GATE 1.83945e-17 
c_425 M30:GATE N_17:2 8.001e-20 
c_426 M30:GATE M32:GATE 1.76894e-19 
c_427 M30:GATE 0 1.76878e-18 
c_428 A M6:SRC 4.28241e-19 
c_429 A M17:BULK 5.44394e-18 
c_430 A GND:1 8.46237e-18 
c_431 A N_17:3 6.75929e-17 
c_432 A M31:DRN 6.30572e-18 
c_433 A N_17:1 8.26192e-18 
c_434 A M6:DRN 2.2527e-19 
c_435 A 0 2.88445e-17 
c_436 M5:GATE M6:SRC 1.09235e-17 
c_437 M5:GATE M8:GATE 3.56175e-18 
c_438 M5:GATE M7:GATE 1.79606e-19 
c_439 M5:GATE M17:BULK 4.31813e-18 
c_440 M5:GATE GND:1 5.29846e-18 
c_441 M5:GATE N_17:3 7.16945e-18 
c_442 M5:GATE N_17:1 1.54098e-17 
c_443 M5:GATE M33:GATE 9.10346e-19 
c_444 M5:GATE N_17:2 1.12749e-19 
c_445 M5:GATE M5:SRC 1.03127e-17 
c_446 M5:GATE M6:DRN 5.03913e-18 
c_447 M5:GATE 0 2.8543e-18 
c_448 M6:GATE GND:1 6.90904e-18 
c_449 M6:GATE M17:BULK 3.37826e-18 
c_450 M6:GATE M8:GATE 2.7447e-19 
c_451 M6:GATE N_17:1 1.09586e-19 
c_452 M6:GATE N_17:3 9.47476e-18 
c_453 M6:GATE M6:SRC 2.23602e-17 
c_454 M6:GATE M5:SRC 1.39309e-18 
c_455 M6:GATE M6:DRN 1.43553e-18 
c_456 N_12:1 M17:GATE 6.54416e-18 
c_457 N_12:1 M8:GATE 1.15619e-20 
c_458 N_12:1 M8:SRC 5.31915e-18 
c_459 N_12:1 M7:GATE 2.7991e-19 
c_460 N_12:1 M16:DRN 3.35273e-17 
c_461 N_12:1 M16:SRC 1.65489e-18 
c_462 N_12:1 M20:SRC 8.95772e-17 
c_463 N_12:1 M17:DRN 1.07261e-17 
c_464 N_12:1 M17:SRC 3.0313e-17 
c_465 N_12:1 M18:DRN 1.09829e-16 
c_466 N_12:1 M4:GATE 3.44137e-18 
c_467 N_12:1 M3:DRN 4.15336e-17 
c_468 N_12:1 M12:GATE 1.19493e-17 
c_469 N_12:1 N_17:3 7.48014e-18 
c_470 N_12:1 M34:GATE 7.11868e-19 
c_471 N_12:1 B 1.01663e-16 
c_472 N_12:1 M23:GATE 1.36592e-17 
c_473 N_12:1 M3:GATE 1.08476e-18 
c_474 N_12:1 M22:DRN 8.37064e-17 
c_475 N_12:1 N_17:1 1.12749e-18 
c_476 N_12:1 N_17:2 9.67386e-19 
c_477 N_12:1 M23:DRN 1.18336e-16 
c_478 N_12:1 M12:SRC 2.78767e-19 
c_479 N_12:1 M20:GATE 7.32251e-18 
c_480 N_12:1 M21:GATE 1.07849e-17 
c_481 N_12:1 M22:GATE 2.75173e-20 
c_482 N_12:1 0 7.99994e-18 
c_483 M34:DRN M17:GATE 1.90874e-21 
c_484 M34:DRN M20:SRC 7.36401e-19 
c_485 M34:DRN M17:SRC 2.15374e-18 
c_486 M34:DRN M18:DRN 3.84439e-17 
c_487 M34:DRN M4:GATE 5.3046e-18 
c_488 M34:DRN M3:DRN 1.61787e-20 
c_489 M34:DRN M34:GATE 1.61047e-17 
c_490 M34:DRN B 2.97839e-17 
c_491 M34:DRN M23:GATE 2.54801e-19 
c_492 M34:DRN M20:DRN 3.90219e-19 
c_493 M34:DRN M23:DRN 9.77278e-19 
c_494 M34:DRN 0 4.496e-18 
c_495 M21:DRN M3:DRN 1.92333e-18 
c_496 M21:DRN M12:GATE 6.90955e-18 
c_497 M21:DRN M34:GATE 2.27491e-20 
c_498 M21:DRN M23:GATE 1.77721e-17 
c_499 M21:DRN M3:GATE 1.47861e-18 
c_500 M21:DRN M22:DRN 3.57352e-17 
c_501 M21:DRN M23:DRN 3.75026e-17 
c_502 M21:DRN M21:GATE 3.08363e-17 
c_503 M21:DRN 0 4.55456e-19 
c_504 M4:DRN M17:GATE 4.99234e-18 
c_505 M4:DRN M16:SRC 3.97884e-21 
c_506 M4:DRN M20:SRC 3.91058e-18 
c_507 M4:DRN M17:DRN 3.94267e-20 
c_508 M4:DRN M17:SRC 3.57351e-17 
c_509 M4:DRN M4:GATE 3.26856e-17 
c_510 M4:DRN M3:DRN 8.74274e-19 
c_511 M4:DRN M34:GATE 1.89772e-20 
c_512 M4:DRN B 2.22858e-19 
c_513 M4:DRN M23:GATE 1.36804e-20 
c_514 M4:DRN 0 1.1223e-17 
c_515 M12:DRN M17:GATE 2.44989e-22 
c_516 M12:DRN M20:SRC 1.26078e-18 
c_517 M12:DRN M4:GATE 4.44668e-21 
c_518 M12:DRN M3:DRN 2.03096e-17 
c_519 M12:DRN M3:GATE 1.4592e-17 
c_520 M12:DRN M22:DRN 2.99112e-18 
c_521 M12:DRN M23:DRN 2.81556e-17 
c_522 M12:DRN M12:SRC 4.90952e-19 
c_523 M12:DRN N_24:1 6.67001e-21 
c_524 M12:DRN M19:GATE 2.26591e-19 
c_525 M12:DRN 0 2.10965e-17 
c_526 M18:GATE M8:SRC 7.88183e-19 
c_527 M18:GATE M20:SRC 2.55455e-17 
c_528 M18:GATE M17:SRC 1.30217e-17 
c_529 M18:GATE M18:DRN 3.86513e-17 
c_530 M18:GATE N_17:3 5.76293e-18 
c_531 M18:GATE M34:GATE 4.68957e-18 
c_532 M18:GATE B 1.227e-18 
c_533 M18:GATE M23:GATE 5.83862e-20 
c_534 M18:GATE N_17:1 3.44575e-19 
c_535 M18:GATE N_17:2 5.24065e-20 
c_536 M18:GATE M32:GATE 7.39067e-20 
c_537 M18:GATE M20:DRN 5.87671e-20 
c_538 M18:GATE M20:GATE 1.04992e-17 
c_539 M18:GATE 0 1.67933e-17 
c_540 M16:GATE M17:GATE 9.10775e-18 
c_541 M16:GATE M8:GATE 1.40206e-19 
c_542 M16:GATE M7:GATE 7.02683e-19 
c_543 M16:GATE M16:DRN 4.67251e-18 
c_544 M16:GATE M16:SRC 1.85206e-17 
c_545 M16:GATE M20:SRC 4.5371e-18 
c_546 M16:GATE M17:SRC 3.11802e-19 
c_547 M16:GATE M18:DRN 1.00484e-17 
c_548 M16:GATE M4:GATE 6.0376e-20 
c_549 M16:GATE N_17:3 2.27423e-18 
c_550 M16:GATE B 1.00078e-17 
c_551 M16:GATE 0 2.89641e-17 
c_552 CI:1 M6:SRC 4.19252e-20 
c_553 CI:1 M7:DRN 1.55738e-19 
c_554 CI:1 M17:BULK 2.05633e-18 
c_555 CI:1 GND:1 3.99839e-20 
c_556 CI:1 M13:SRC 2.39646e-18 
c_557 CI:1 0 6.64685e-18 
c_558 M27:GATE 0 1.48856e-17 
c_559 M26:GATE 0 2.81691e-17 
c_560 CI M7:DRN 2.58052e-19 
c_561 CI M17:BULK 4.2609e-18 
c_562 CI GND:1 1.09232e-18 
c_563 CI M13:SRC 8.49344e-19 
c_564 CI M14:DRN 3.87544e-18 
c_565 CI M2:DRN 4.23738e-22 
c_566 CI 0 7.81032e-18 
c_567 M14:GATE M6:SRC 4.35819e-18 
c_568 M14:GATE M7:DRN 1.03554e-17 
c_569 M14:GATE M17:BULK 4.51844e-18 
c_570 M14:GATE GND:1 4.57161e-18 
c_571 M14:GATE M13:SRC 9.56924e-19 
c_572 M14:GATE M14:DRN 1.17652e-17 
c_573 M14:GATE 0 7.77083e-18 
c_574 M15:GATE GND:1 5.52198e-18 
c_575 M15:GATE M17:BULK 2.59274e-18 
c_576 M15:GATE M14:DRN 8.19982e-19 
c_577 M15:GATE M13:SRC 1.03192e-17 
c_578 M15:GATE M6:SRC 4.35819e-18 
c_579 M15:GATE M7:DRN 5.66455e-18 
c_580 M15:GATE 0 4.87576e-19 
c_581 N_5:1 M6:SRC 1.87047e-19 
c_582 N_5:1 M7:DRN 3.90261e-18 
c_583 N_5:1 M20:SRC 5.9789e-18 
c_584 N_5:1 M17:BULK 1.28876e-17 
c_585 N_5:1 M12:GATE 3.42179e-19 
c_586 N_5:1 GND:1 1.0793e-16 
c_587 N_5:1 M22:DRN 8.31645e-19 
c_588 N_5:1 M23:DRN 5.6845e-19 
c_589 N_5:1 M12:SRC 1.3618e-16 
c_590 N_5:1 N_24:1 5.3523e-18 
c_591 N_5:1 M24:GATE 1.52819e-17 
c_592 N_5:1 M25:DRN 5.38834e-17 
c_593 N_5:1 M19:GATE 1.54506e-17 
c_594 N_5:1 M11:GATE 9.39716e-18 
c_595 N_5:1 N_20:1 2.46268e-16 
c_596 N_5:1 M11:DRN 5.46293e-18 
c_597 N_5:1 M24:DRN 5.90049e-19 
c_598 N_5:1 M9:GATE 1.64495e-17 
c_599 N_5:1 M13:DRN 9.44505e-17 
c_600 N_5:1 M13:SRC 4.70488e-18 
c_601 N_5:1 CI:1 2.42753e-17 
c_602 N_5:1 M15:GATE 2.74514e-18 
c_603 N_5:1 CI 1.37759e-16 
c_604 N_5:1 M14:GATE 4.96474e-18 
c_605 N_5:1 M14:DRN 1.0944e-17 
c_606 N_5:1 M28:GATE 1.65507e-20 
c_607 N_5:1 M9:SRC 2.55915e-18 
c_608 N_5:1 M27:GATE 5.65534e-18 
c_609 N_5:1 M26:GATE 6.32399e-18 
c_610 N_5:1 M10:GATE 4.73749e-18 
c_611 N_5:1 M22:GATE 4.69715e-18 
c_612 N_5:1 0 3.37008e-18 
c_613 M25:GATE GND:1 1.09499e-19 
c_614 M25:GATE M23:GATE 6.21428e-21 
c_615 M25:GATE M12:SRC 5.13316e-18 
c_616 M25:GATE M24:GATE 8.08876e-18 
c_617 M25:GATE M25:DRN 1.6976e-17 
c_618 M25:GATE M19:GATE 1.356e-19 
c_619 M25:GATE N_20:1 8.27511e-18 
c_620 M25:GATE M24:DRN 6.04472e-20 
c_621 M25:GATE M13:DRN 3.0166e-18 
c_622 M25:GATE CI:1 9.88872e-18 
c_623 M25:GATE CI 2.23164e-18 
c_624 M25:GATE CO 3.1233e-19 
c_625 M25:GATE M28:GATE 4.34339e-20 
c_626 M25:GATE M27:GATE 9.26251e-18 
c_627 M25:GATE M26:GATE 1.99087e-19 
c_628 M25:GATE M22:GATE 2.6233e-18 
c_629 M25:GATE 0 3.61596e-18 
c_630 M22:SRC M6:SRC 6.04654e-20 
c_631 M22:SRC GND:1 2.3551e-17 
c_632 M22:SRC M3:GATE 2.67223e-22 
c_633 M22:SRC M22:DRN 3.75286e-18 
c_634 M22:SRC M23:DRN 3.34465e-21 
c_635 M22:SRC M24:GATE 1.5013e-17 
c_636 M22:SRC M25:DRN 5.78741e-20 
c_637 M22:SRC M19:GATE 3.36487e-17 
c_638 M22:SRC N_20:1 8.27162e-19 
c_639 M22:SRC M24:DRN 6.82019e-18 
c_640 M22:SRC CO 3.12578e-17 
c_641 M22:SRC M1:DRN 3.32368e-18 
c_642 M22:SRC M1:GATE 1.36319e-18 
c_643 M22:SRC M28:GATE 2.95668e-19 
c_644 M22:SRC M28:DRN 1.25917e-18 
c_645 M22:SRC M21:GATE 1.2593e-20 
c_646 M22:SRC M29:GATE 7.14144e-19 
c_647 M22:SRC M22:GATE 1.66312e-17 
c_648 M22:SRC 0 1.27841e-17 
c_649 M27:SRC M6:SRC 6.09174e-20 
c_650 M27:SRC M7:DRN 2.61021e-23 
c_651 M27:SRC M12:SRC 5.06563e-18 
c_652 M27:SRC M25:DRN 5.7874e-20 
c_653 M27:SRC N_20:1 5.54893e-18 
c_654 M27:SRC M11:DRN 1.2939e-19 
c_655 M27:SRC CI:1 1.42804e-17 
c_656 M27:SRC CI 1.19979e-18 
c_657 M27:SRC CO 1.16008e-19 
c_658 M27:SRC M28:DRN 8.01198e-20 
c_659 M27:SRC M27:GATE 1.8805e-17 
c_660 M27:SRC M26:GATE 1.67205e-17 
c_661 M14:SRC M6:SRC 9.88896e-18 
c_662 M14:SRC M7:DRN 9.75593e-19 
c_663 M14:SRC GND:1 2.70002e-17 
c_664 M14:SRC M13:DRN 8.68111e-21 
c_665 M14:SRC CI:1 3.3125e-17 
c_666 M14:SRC M15:GATE 7.14116e-18 
c_667 M14:SRC CI 1.38674e-17 
c_668 M14:SRC CO 2.028e-17 
c_669 M14:SRC M1:DRN 6.7306e-20 
c_670 M14:SRC M9:SRC 3.47244e-20 
c_671 M13:GATE M6:SRC 4.35747e-18 
c_672 M13:GATE M7:DRN 5.08342e-18 
c_673 M13:GATE M17:BULK 5.20935e-18 
c_674 M13:GATE GND:1 2.08261e-18 
c_675 M13:GATE M3:GATE 2.71183e-18 
c_676 M13:GATE N_24:1 2.7724e-18 
c_677 M13:GATE M25:DRN 1.65965e-19 
c_678 M13:GATE M13:DRN 1.06502e-17 
c_679 M13:GATE M13:SRC 1.27385e-17 
c_680 M13:GATE CI:1 1.81494e-17 
c_681 M13:GATE M15:GATE 3.68959e-18 
c_682 M13:GATE CI 4.51085e-19 
c_683 M13:GATE M14:GATE 2.05377e-19 
c_684 M13:GATE 0 1.6146e-20 
c_685 M11:SRC M6:SRC 7.7101e-18 
c_686 M11:SRC M7:DRN 3.09322e-20 
c_687 M11:SRC M3:DRN 8.55352e-20 
c_688 M11:SRC GND:1 3.60668e-17 
c_689 M11:SRC M3:GATE 1.47472e-17 
c_690 M11:SRC M22:DRN 4.68127e-19 
c_691 M11:SRC M12:SRC 2.8948e-19 
c_692 M11:SRC M24:GATE 1.27568e-17 
c_693 M11:SRC M11:GATE 6.83343e-18 
c_694 M11:SRC N_20:1 6.16294e-19 
c_695 M11:SRC M11:DRN 5.67668e-18 
c_696 M11:SRC M24:DRN 2.18011e-19 
c_697 M11:SRC M9:GATE 5.28306e-19 
c_698 M11:SRC M13:SRC 4.11909e-22 
c_699 M11:SRC CO 3.94173e-17 
c_700 M11:SRC M9:SRC 9.39431e-20 
c_701 M11:SRC M10:GATE 2.62844e-17 
c_702 M11:SRC 0 1.30669e-19 
c_703 VDD:1 M17:SRC 1.6275e-20 
c_704 VDD:1 M12:SRC 5.7831e-18 
c_705 VDD:1 N_20:1 3.08062e-18 
c_706 VDD:1 M28:GATE 5.5668e-19 
c_707 VDD:1 M27:GATE 1.05048e-18 
c_708 VDD:1 M26:GATE 5.69846e-19 
c_709 VDD:1 M29:GATE 4.29317e-19 
c_710 VDD:1 0 2.27362e-17 
c_711 VDD:2 N_12:1 1.6275e-20 
c_712 VDD:2 M18:GATE 5.78259e-20 
c_713 VDD:2 M34:GATE 2.06076e-18 
c_714 VDD:2 M23:GATE 7.17426e-19 
c_715 VDD:2 M3:GATE 3.15476e-19 
c_716 VDD:2 M30:GATE 4.50706e-19 
c_717 VDD:2 M33:GATE 8.27763e-19 
c_718 VDD:2 M32:GATE 9.45141e-19 
c_719 VDD:2 M12:SRC 4.54134e-17 
c_720 VDD:2 M24:GATE 1.13644e-18 
c_721 VDD:2 N_20:1 3.69677e-17 
c_722 VDD:2 CO 4.87715e-19 
c_723 VDD:2 M28:GATE 1.25791e-17 
c_724 VDD:2 S 1.19354e-17 
c_725 VDD:2 M31:GATE 5.20601e-19 
c_726 VDD:2 M25:GATE 1.34083e-18 
c_727 VDD:2 M27:GATE 4.02369e-19 
c_728 VDD:2 M26:GATE 5.86619e-19 
c_729 VDD:2 M29:GATE 2.38698e-18 
c_730 VDD:2 0 1.08673e-18 
c_731 M34:BULK M20:SRC 2.80964e-18 
c_732 M34:BULK M17:SRC 8.76826e-18 
c_733 M34:BULK M18:DRN 2.62343e-18 
c_734 M34:BULK N_12:1 8.93837e-18 
c_735 M34:BULK M34:DRN 1.72081e-18 
c_736 M34:BULK M4:GATE 4.14774e-18 
c_737 M34:BULK M3:DRN 5.43458e-18 
c_738 M34:BULK M12:GATE 6.64669e-18 
c_739 M34:BULK N_17:3 8.6526e-18 
c_740 M34:BULK M34:GATE 8.61385e-18 
c_741 M34:BULK B 3.81313e-18 
c_742 M34:BULK M23:GATE 1.61922e-17 
c_743 M34:BULK M22:DRN 1.09557e-17 
c_744 M34:BULK M31:DRN 3.01576e-18 
c_745 M34:BULK M30:GATE 7.33713e-18 
c_746 M34:BULK N_17:1 2.31208e-18 
c_747 M34:BULK M33:GATE 3.86672e-18 
c_748 M34:BULK N_17:2 2.03475e-18 
c_749 M34:BULK M32:GATE 1.50672e-18 
c_750 M34:BULK M20:DRN 2.05409e-18 
c_751 M34:BULK M23:DRN 4.45702e-19 
c_752 M34:BULK M24:GATE 3.62281e-18 
c_753 M34:BULK A 6.08178e-18 
c_754 M34:BULK A:1 6.77599e-18 
c_755 M34:BULK M20:GATE 3.78941e-18 
c_756 M34:BULK M19:GATE 1.43863e-18 
c_757 M34:BULK N_20:1 1.78568e-17 
c_758 M34:BULK M24:DRN 1.31912e-18 
c_759 M34:BULK CI:1 8.21664e-18 
c_760 M34:BULK CI 1.58157e-18 
c_761 M34:BULK N_5:1 7.03078e-18 
c_762 M34:BULK CO 3.273e-18 
c_763 M34:BULK M28:GATE 8.36534e-18 
c_764 M34:BULK S 7.074e-18 
c_765 M34:BULK M21:DRN 8.73867e-19 
c_766 M34:BULK M22:SRC 7.82637e-19 
c_767 M34:BULK M29:SRC 2.99859e-18 
c_768 M34:BULK M31:GATE 4.05763e-18 
c_769 M34:BULK M21:GATE 1.48829e-18 
c_770 M34:BULK M25:GATE 4.43849e-18 
c_771 M34:BULK M27:GATE 2.57651e-18 
c_772 M34:BULK M26:GATE 3.26115e-18 
c_773 M34:BULK M29:GATE 1.80696e-18 
c_774 M34:BULK M22:GATE 2.8416e-18 
c_775 M34:SRC M16:SRC 3.6903e-19 
c_776 M34:SRC M20:SRC 3.64945e-21 
c_777 M34:SRC M18:DRN 4.26821e-20 
c_778 M34:SRC N_12:1 5.61452e-18 
c_779 M34:SRC M4:GATE 4.95328e-18 
c_780 M34:SRC M3:DRN 2.05347e-19 
c_781 M34:SRC M12:GATE 1.03099e-20 
c_782 M34:SRC M34:GATE 1.23062e-17 
c_783 M34:SRC B 3.62433e-18 
c_784 M34:SRC M23:GATE 1.16335e-17 
c_785 M34:SRC M3:GATE 9.0219e-24 
c_786 M34:SRC M22:DRN 2.54646e-17 
c_787 M34:SRC M23:DRN 2.36051e-20 
c_788 M34:SRC M24:GATE 2.48829e-17 
c_789 M34:SRC M20:GATE 9.13425e-19 
c_790 M34:SRC M19:GATE 1.41607e-19 
c_791 M34:SRC N_20:1 2.25125e-18 
c_792 M34:SRC M11:DRN 3.63324e-20 
c_793 M34:SRC M24:DRN 1.76941e-20 
c_794 M34:SRC M9:GATE 3.54152e-21 
c_795 M34:SRC CI:1 6.42359e-20 
c_796 M34:SRC M27:SRC 1.26752e-19 
c_797 M34:SRC N_5:1 3.80409e-20 
c_798 M34:SRC M14:SRC 1.50365e-24 
c_799 M34:SRC S 8.52885e-19 
c_800 M34:SRC M21:DRN 1.39761e-19 
c_801 M34:SRC M22:SRC 1.78842e-20 
c_802 M34:SRC M28:DRN 1.14489e-20 
c_803 M34:SRC M21:GATE 3.61813e-17 
c_804 M34:SRC M25:GATE 4.45432e-18 
c_805 M34:SRC M27:GATE 5.1394e-18 
c_806 M34:SRC M26:GATE 5.1411e-18 
c_807 M34:SRC M29:GATE 5.1415e-18 
c_808 M34:SRC M22:GATE 1.32285e-17 
c_809 M34:SRC 0 2.6556e-17 
c_810 M25:SRC N_17:3 6.26951e-20 
c_811 M25:SRC M34:GATE 1.46697e-20 
c_812 M25:SRC M12:SRC 5.87379e-18 
c_813 M25:SRC M24:GATE 1.70299e-18 
c_814 M25:SRC M20:GATE 2.84372e-20 
c_815 M25:SRC N_20:1 6.27263e-18 
c_816 M25:SRC M24:DRN 1.80461e-19 
c_817 M25:SRC CI 1.95259e-19 
c_818 M25:SRC N_5:1 1.4896e-17 
c_819 M25:SRC S 1.72459e-20 
c_820 M25:SRC M25:GATE 1.99345e-17 
c_821 M25:SRC M27:GATE 2.0888e-17 
c_822 M25:SRC M26:GATE 1.06003e-18 
c_823 M25:SRC 0 4.7093e-18 
c_824 M28:SRC N_17:3 6.82198e-20 
c_825 M28:SRC M28:GATE 3.10677e-17 
c_826 M28:SRC M29:GATE 2.85465e-17 
c_827 M28:SRC N_20:1 1.34875e-17 
c_828 M28:SRC S 2.67493e-19 
c_829 M28:SRC CO 1.63206e-19 
c_830 M28:SRC 0 3.49552e-18 
c_831 M26:DRN M12:SRC 1.65101e-17 
c_832 M26:DRN N_20:1 2.49403e-18 
c_833 M26:DRN CI:1 1.78234e-18 
c_834 M26:DRN CI 1.41453e-19 
c_835 M26:DRN N_5:1 2.44763e-18 
c_836 M26:DRN M28:GATE 1.35689e-17 
c_837 M26:DRN M28:DRN 2.28256e-17 
c_838 M26:DRN M27:GATE 1.3449e-18 
c_839 M26:DRN M26:GATE 1.27644e-17 
c_840 M26:DRN 0 3.14005e-18 
c_841 VDD M16:DRN 3.32634e-18 
c_842 VDD M16:SRC 1.85758e-18 
c_843 VDD M20:SRC 1.13344e-18 
c_844 VDD M18:DRN 1.49645e-18 
c_845 VDD N_12:1 1.14307e-16 
c_846 VDD M34:DRN 1.63272e-18 
c_847 VDD M3:DRN 1.55775e-18 
c_848 VDD N_17:3 1.97622e-16 
c_849 VDD M18:GATE 1.30777e-18 
c_850 VDD M34:GATE 3.63266e-17 
c_851 VDD B 2.99622e-18 
c_852 VDD M23:GATE 2.64344e-17 
c_853 VDD M22:DRN 2.06523e-16 
c_854 VDD M31:DRN 1.78593e-18 
c_855 VDD M30:GATE 7.51124e-18 
c_856 VDD M33:GATE 7.10788e-18 
c_857 VDD M32:GATE 8.04995e-18 
c_858 VDD M20:DRN 1.05994e-18 
c_859 VDD M23:DRN 9.07078e-19 
c_860 VDD M24:GATE 2.60846e-17 
c_861 VDD A 8.5028e-18 
c_862 VDD A:1 7.33255e-19 
c_863 VDD M32:SRC 1.43737e-18 
c_864 VDD M20:GATE 4.56927e-18 
c_865 VDD M19:GATE 1.26734e-18 
c_866 VDD N_20:1 1.14113e-17 
c_867 VDD M24:DRN 9.88827e-19 
c_868 VDD M27:SRC 1.65063e-19 
c_869 VDD N_5:1 1.38742e-18 
c_870 VDD CO 4.35303e-19 
c_871 VDD M28:GATE 1.81076e-17 
c_872 VDD S 2.74994e-17 
c_873 VDD M21:DRN 1.71257e-18 
c_874 VDD M22:SRC 9.35496e-19 
c_875 VDD M28:DRN 4.04442e-19 
c_876 VDD M29:SRC 1.96268e-18 
c_877 VDD M31:GATE 8.77035e-18 
c_878 VDD M21:GATE 3.70682e-18 
c_879 VDD M25:GATE 4.62128e-18 
c_880 VDD M27:GATE 3.92852e-18 
c_881 VDD M26:GATE 5.90685e-18 
c_882 VDD M29:GATE 8.84597e-18 
c_883 VDD M22:GATE 2.98147e-18 
c_884 VDD 0 2.1568e-16 
c_885 M31:SRC M8:SRC 3.81007e-20 
c_886 M31:SRC M16:DRN 9.80801e-19 
c_887 M31:SRC M20:SRC 6.12588e-18 
c_888 M31:SRC M17:SRC 3.80228e-20 
c_889 M31:SRC M18:DRN 4.13827e-18 
c_890 M31:SRC N_12:1 1.31629e-19 
c_891 M31:SRC M34:DRN 7.51162e-18 
c_892 M31:SRC M4:DRN 2.87683e-20 
c_893 M31:SRC M3:DRN 1.65313e-19 
c_894 M31:SRC M12:DRN 6.98307e-20 
c_895 M31:SRC M12:GATE 2.20026e-20 
c_896 M31:SRC N_17:3 3.59397e-18 
c_897 M31:SRC M18:GATE 1.64483e-18 
c_898 M31:SRC M34:GATE 3.90184e-17 
c_899 M31:SRC B 5.48497e-20 
c_900 M31:SRC M23:GATE 2.90751e-17 
c_901 M31:SRC M22:DRN 1.01457e-17 
c_902 M31:SRC M31:DRN 9.62578e-18 
c_903 M31:SRC M30:GATE 1.09595e-17 
c_904 M31:SRC N_17:1 2.36517e-20 
c_905 M31:SRC M33:GATE 9.49908e-18 
c_906 M31:SRC M32:GATE 9.11608e-18 
c_907 M31:SRC M20:DRN 7.79196e-18 
c_908 M31:SRC M23:DRN 6.05163e-18 
c_909 M31:SRC M12:SRC 1.21789e-19 
c_910 M31:SRC M24:GATE 2.72289e-17 
c_911 M31:SRC A 2.49136e-18 
c_912 M31:SRC A:1 8.43637e-18 
c_913 M31:SRC M32:SRC 8.52245e-18 
c_914 M31:SRC M6:DRN 3.81007e-20 
c_915 M31:SRC M19:GATE 1.57042e-18 
c_916 M31:SRC M11:SRC 9.90438e-20 
c_917 M31:SRC N_20:1 3.65664e-21 
c_918 M31:SRC M11:DRN 3.96861e-20 
c_919 M31:SRC M24:DRN 5.75503e-18 
c_920 M31:SRC CI:1 4.02231e-20 
c_921 M31:SRC M27:SRC 5.41074e-18 
c_922 M31:SRC N_5:1 2.0189e-20 
c_923 M31:SRC M14:SRC 6.14111e-20 
c_924 M31:SRC M1:DRN 3.91388e-21 
c_925 M31:SRC M28:GATE 1.91051e-17 
c_926 M31:SRC M2:SRC 3.06117e-20 
c_927 M31:SRC S 9.04336e-20 
c_928 M31:SRC M21:DRN 7.50253e-18 
c_929 M31:SRC M22:SRC 5.68889e-18 
c_930 M31:SRC M28:DRN 2.77148e-18 
c_931 M31:SRC M29:SRC 9.72802e-18 
c_932 M31:SRC M31:GATE 2.23713e-17 
c_933 M31:SRC M25:GATE 4.82349e-18 
c_934 M31:SRC M27:GATE 4.35783e-18 
c_935 M31:SRC M26:GATE 4.35783e-18 
c_936 M31:SRC M29:GATE 4.35799e-18 
c_937 M31:SRC 0 1.8626e-16 
c_938 M30:SRC M34:GATE 9.25068e-20 
c_939 M30:SRC N_17:3 9.99436e-18 
c_940 M30:SRC M31:GATE 8.3293e-19 
c_941 M30:SRC M30:GATE 1.03177e-17 
c_942 M30:SRC M33:GATE 1.03177e-17 
c_943 M30:SRC M32:GATE 8.3293e-19 
c_944 M30:SRC M16:DRN 2.22637e-19 
c_945 M30:SRC 0 4.45698e-18 
c_946 M32:DRN M8:SRC 7.1264e-18 
c_947 M32:DRN M16:DRN 5.26444e-22 
c_948 M32:DRN M20:SRC 3.00347e-19 
c_949 M32:DRN M18:DRN 1.23195e-19 
c_950 M32:DRN N_12:1 3.5278e-19 
c_951 M32:DRN M34:DRN 8.04316e-20 
c_952 M32:DRN M4:DRN 1.50365e-24 
c_953 M32:DRN N_17:3 5.31231e-18 
c_954 M32:DRN M18:GATE 1.70646e-19 
c_955 M32:DRN M34:GATE 3.16264e-17 
c_956 M32:DRN M33:GATE 8.3293e-19 
c_957 M32:DRN M32:GATE 1.36897e-17 
c_958 M32:DRN M20:DRN 3.73953e-17 
c_959 M32:DRN M20:GATE 3.17435e-17 
c_960 M32:DRN 0 7.2922e-18 

.ENDS
