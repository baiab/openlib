
.subckt DFD4  D CP Q QN
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=2.358e-06 sb=8.1e-07 w=0.54u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=2.034e-06 sb=1.134e-06 w=0.54u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK nch ad=0.06966p as=0.1134p l=0.09u nrd=0.24 nrs=0.387 pd=0.9108u ps=1.539u sa=4.095e-07 sb=2.403e-07 w=0.54u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK nch ad=0.06075p as=0.11016p l=0.09u nrd=0.209 nrs=0.379 pd=0.927u ps=1.494u sa=4.86e-07 sb=2.043e-07 w=0.54u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK nch ad=0.0162p as=0.04536p l=0.09u nrd=0.5 nrs=1.389 pd=0.36u ps=0.6849u sa=9.9e-07 sb=1.6164e-06 w=0.18u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK nch ad=0.08424p as=0.06642p l=0.09u nrd=0.511 nrs=0.405 pd=1.224u ps=1.026u sa=7.929e-07 sb=2.07e-07 w=0.405u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK nch ad=0.04617p as=0.08829p l=0.09u nrd=0.205 nrs=0.388 pd=0.684u ps=1.638u sa=1.44e-07 sb=6.03e-07 w=0.477u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.06318p as=0.15714p l=0.09u nrd=0.217 nrs=0.539 pd=0.774u ps=1.926u sa=2.25e-07 sb=2.943e-06 w=0.54u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=1.431e-06 sb=1.737e-06 w=0.54u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=8.28e-07 sb=2.34e-06 w=0.54u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=2.637e-06 sb=5.31e-07 w=0.54u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.0243p as=0.0162p l=0.09u nrd=0.756 nrs=0.5 pd=0.3915u ps=0.36u sa=7.155e-07 sb=1.9125e-06 w=0.18u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK nch ad=0.11178p as=0.06075p l=0.09u nrd=0.383 nrs=0.209 pd=1.494u ps=0.927u sa=2.07e-07 sb=4.833e-07 w=0.54u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK nch ad=0.07371p as=0.05265p l=0.09u nrd=0.252 nrs=0.181 pd=1.1745u ps=0.774u sa=3.546e-07 sb=2.349e-07 w=0.54u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK nch ad=0.04941p as=0.09477p l=0.09u nrd=0.343 nrs=0.661 pd=0.6372u ps=1.4391u sa=2.745e-07 sb=7.812e-07 w=0.378u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK nch ad=0.06642p as=0.06399p l=0.09u nrd=0.405 nrs=0.388 pd=1.026u ps=0.9099u sa=3.69e-07 sb=5.04e-07 w=0.405u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=5.49e-07 sb=2.619e-06 w=0.54u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK nch ad=0.02835p as=0.03807p l=0.09u nrd=0.873 nrs=1.163 pd=0.4041u ps=0.513u sa=1.7118e-06 sb=8.46e-07 w=0.18u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=1.755e-06 sb=1.413e-06 w=0.54u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=1.152e-06 sb=2.016e-06 w=0.54u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.11178p as=0.06318p l=0.09u nrd=0.383 nrs=0.217 pd=1.494u ps=0.774u sa=2.961e-06 sb=2.07e-07 w=0.54u 
MM37 M37:DRN M37:GATE M37:SRC M37:BULK pch ad=0.14904p as=0.08424p l=0.09u nrd=0.287 nrs=0.162 pd=1.854u ps=0.954u sa=2.961e-06 sb=2.07e-07 w=0.72u 
MM39 M39:DRN M39:GATE M39:SRC M39:BULK pch ad=0.07776p as=0.08424p l=0.09u nrd=0.15 nrs=0.162 pd=1.107u ps=0.954u sa=2.358e-06 sb=8.1e-07 w=0.72u 
MM30 M30:DRN M30:GATE M30:SRC M30:BULK pch ad=0.08262p as=0.06804p l=0.09u nrd=0.283 nrs=0.233 pd=1.0557u ps=0.954u sa=4.05e-07 sb=5.04e-07 w=0.54u 
MM23 M23:DRN M23:GATE M23:SRC M23:BULK pch ad=0.0243p as=0.04536p l=0.09u nrd=0.333 nrs=0.617 pd=0.45u ps=0.5463u sa=1.053e-06 sb=1.503e-06 w=0.27u 
MM32 M32:DRN M32:GATE M32:SRC M32:BULK pch ad=0.08424p as=0.19764p l=0.09u nrd=0.162 nrs=0.381 pd=0.954u ps=2.286u sa=2.25e-07 sb=2.943e-06 w=0.72u 
MM25 M25:DRN M25:GATE M25:SRC M25:BULK pch ad=0.04455p as=0.13122p l=0.09u nrd=0.212 nrs=0.625 pd=0.6633u ps=1.944u sa=1.8e-07 sb=9.18e-07 w=0.459u 
MM41 M41:DRN M41:GATE M41:SRC M41:BULK pch ad=0.14904p as=0.07776p l=0.09u nrd=0.287 nrs=0.15 pd=1.854u ps=1.107u sa=2.07e-07 sb=4.752e-07 w=0.72u 
MM34 M34:DRN M34:GATE M34:SRC M34:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=1.431e-06 sb=1.737e-06 w=0.72u 
MM27 M27:DRN M27:GATE M27:SRC M27:BULK pch ad=0.05103p as=0.04131p l=0.09u nrd=0.705 nrs=0.567 pd=0.5832u ps=0.5283u sa=1.6569e-06 sb=8.46e-07 w=0.27u 
MM36 M36:DRN M36:GATE M36:SRC M36:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=8.28e-07 sb=2.34e-06 w=0.72u 
MM29 M29:DRN M29:GATE M29:SRC M29:BULK pch ad=0.11178p as=0.06804p l=0.09u nrd=0.383 nrs=0.233 pd=1.494u ps=0.954u sa=8.487e-07 sb=2.07e-07 w=0.54u 
MM38 M38:DRN M38:GATE M38:SRC M38:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=2.637e-06 sb=5.31e-07 w=0.72u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK pch ad=0.0243p as=0.03726p l=0.09u nrd=0.333 nrs=0.516 pd=0.45u ps=0.5148u sa=7.83e-07 sb=1.8063e-06 w=0.27u 
MM31 M31:DRN M31:GATE M31:SRC M31:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=5.49e-07 sb=2.619e-06 w=0.72u 
MM24 M24:DRN M24:GATE M24:SRC M24:BULK pch ad=0.07128p as=0.05022p l=0.09u nrd=0.272 nrs=0.19 pd=0.9792u ps=0.7407u sa=3.834e-07 sb=3.969e-07 w=0.513u 
MM40 M40:DRN M40:GATE M40:SRC M40:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=2.034e-06 sb=1.134e-06 w=0.72u 
MM33 M33:DRN M33:GATE M33:SRC M33:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=1.755e-06 sb=1.413e-06 w=0.72u 
MM26 M26:DRN M26:GATE M26:SRC M26:BULK pch ad=0.081p as=0.06156p l=0.09u nrd=0.343 nrs=0.261 pd=0.9837u ps=0.7542u sa=4.626e-07 sb=8.577e-07 w=0.486u 
MM42 M42:DRN M42:GATE M42:SRC M42:BULK pch ad=0.07776p as=0.14418p l=0.09u nrd=0.15 nrs=0.278 pd=1.107u ps=1.908u sa=4.86e-07 sb=1.917e-07 w=0.72u 
MM35 M35:DRN M35:GATE M35:SRC M35:BULK pch ad=0.07776p as=0.08424p l=0.09u nrd=0.15 nrs=0.162 pd=1.107u ps=0.954u sa=1.152e-06 sb=2.016e-06 w=0.72u 
MM28 M28:DRN M28:GATE M28:SRC M28:BULK pch ad=0.081p as=0.1215p l=0.09u nrd=0.198 nrs=0.298 pd=0.9918u ps=1.3788u sa=5.049e-07 sb=3.528e-07 w=0.639u 
R1 M13:SRC M18:DRN 0.001
R2 M14:DRN M11:SRC 0.001
R3 M23:DRN M22:DRN 0.001
R4 M26:GATE M13:DRN 207.453
R5 M26:GATE M15:GATE 165.48
R6 M26:GATE M24:DRN 203.484
R7 M24:DRN M13:DRN 46.3045
R8 M24:DRN M15:GATE 170.233
R9 M24:DRN M22:SRC 0.001
R10 M15:GATE M13:DRN 173.553
R11 M13:DRN M11:DRN 0.001
R12 M24:GATE M13:GATE 262.602
R13 M24:GATE D 78.4552
R14 D M13:GATE 80.9623
R15 M25:DRN M24:SRC 0.001
R16 M41:GATE M20:GATE 280.312
R17 M41:GATE CP 90.6679
R18 CP M20:GATE 73.5411
R19 M28:DRN M14:GATE 152.931
R20 M28:DRN M23:GATE 239.914
R21 M28:DRN M15:DRN 46.2068
R22 M28:DRN M26:SRC 0.001
R23 M15:DRN M14:GATE 145.875
R24 M15:DRN M23:GATE 228.845
R25 M15:DRN M12:DRN 1.32479e-09
R26 M23:GATE M14:GATE 161.927
R27 Q M36:DRN 9.40096
R28 Q M5:SRC 18.2207
R29 Q M34:DRN 9.27773
R30 Q M3:DRN 18.1503
R31 M36:DRN M34:DRN 605.309
R32 M36:DRN M35:SRC 0.001
R33 M34:DRN M33:DRN 0.001
R34 M3:DRN M4:DRN 0.001
R35 M5:SRC M6:DRN 0.001
R36 QN M10:DRN 9.31167
R37 QN M40:DRN 9.4078
R38 QN M8:DRN 9.23691
R39 QN M38:DRN 9.27763
R40 M40:DRN M38:DRN 605.749
R41 M40:DRN M39:SRC 0.001
R42 M38:DRN M37:SRC 0.001
R43 M10:DRN M8:DRN 704.668
R44 M10:DRN M9:SRC 0.001
R45 M8:DRN M7:SRC 0.001
R46 M21:BULK M20:SRC 7.31417e-06
R47 M21:BULK M7:BULK 0.001
R48 M21:BULK M4:BULK 0.001
R49 M21:BULK M3:BULK 0.001
R50 M21:BULK M10:BULK 0.001
R51 M21:BULK M9:BULK 0.001
R52 M21:BULK M20:BULK 0.001
R53 M21:BULK M18:BULK 0.001
R54 M21:BULK M13:BULK 0.001
R55 M21:BULK M11:BULK 0.001
R56 M21:BULK M14:BULK 0.001
R57 M21:BULK M15:BULK 0.001
R58 M21:BULK M12:BULK 0.001
R59 M21:BULK M19:BULK 0.001
R60 M21:BULK M17:BULK 0.001
R61 M21:BULK M16:BULK 0.001
R62 M21:BULK M2:BULK 0.001
R63 M21:BULK M1:BULK 0.001
R64 M21:BULK M6:BULK 0.001
R65 M21:BULK M5:BULK 0.001
R66 M21:BULK M8:BULK 0.001
R67 M9:DRN M8:SRC 0.001
R68 M9:DRN M20:SRC 1.42857e-09
R69 M3:SRC M10:SRC 0.001
R70 M3:SRC M20:SRC 1.42857e-09
R71 M5:DRN M4:SRC 0.001
R72 M5:DRN M20:SRC 1.42857e-09
R73 M1:SRC M6:SRC 0.001
R74 M1:SRC M20:SRC 1.42857e-09
R75 GND:1 M15:SRC 30.4354
R76 GND:1 M20:SRC 1.35545
R77 GND:1 GND 1.73735
R78 GND:1 M7:DRN 9.28955
R79 GND M20:SRC 1.4132
R80 M16:SRC M17:DRN 0.001
R81 M16:SRC M20:SRC 1.55338e-10
R82 M2:SRC M20:SRC 1.44e-09
R83 M20:SRC M15:SRC 0.001
R84 M20:SRC M18:SRC 1.08081e-09
R85 M20:SRC M21:DRN 0.001
R86 M14:SRC M15:SRC 7.72222e-10
R87 N_28:1 M18:GATE 145.997
R88 N_28:1 M20:DRN 18.3631
R89 N_28:1 M21:GATE 83.2161
R90 N_28:1 M42:GATE 104.899
R91 N_28:1 M41:DRN 18.6145
R92 M22:GATE M28:GATE 280.375
R93 M22:GATE M42:GATE 340.13
R94 M42:GATE M18:GATE 575.605
R95 M42:GATE M28:GATE 956.278
R96 M42:GATE M21:GATE 328.086
R97 M28:GATE M19:GATE 135.6
R98 M21:GATE M18:GATE 456.624
R99 N_26:1 M11:GATE 39.9382
R100 N_26:1 M12:GATE 119.667
R101 N_26:1 M21:SRC 10.9233
R102 N_26:1 M25:GATE 63.9088
R103 N_26:1 M42:SRC 11.2166
R104 N_26:1 M27:GATE 48.4624
R105 M27:GATE M12:GATE 4967.44
R106 M42:SRC M21:SRC 144.923
R107 M42:SRC M25:GATE 847.901
R108 M25:GATE M21:SRC 825.729
R109 VDD:1 M41:SRC 0.932338
R110 VDD:1 M26:DRN 18.3596
R111 VDD:1 M25:SRC 18.2241
R112 VDD:1 M32:SRC 38.2295
R113 VDD:1 M37:DRN 15.662
R114 VDD:1 VDD 0.385643
R115 M42:BULK M41:SRC 7.33998e-06
R116 M42:BULK M30:SRC 0.00474834
R117 M42:BULK M32:SRC 0.00308642
R118 M42:BULK M31:SRC 0.00561167
R119 M42:BULK M35:DRN 0.00561167
R120 M42:BULK M33:SRC 0.00561167
R121 M42:BULK M39:DRN 0.00561167
R122 M42:BULK M41:BULK 0.001
R123 M42:BULK M25:BULK 0.001
R124 M42:BULK M24:BULK 0.001
R125 M42:BULK M22:BULK 0.001
R126 M42:BULK M23:BULK 0.001
R127 M42:BULK M26:BULK 0.001
R128 M42:BULK M28:BULK 0.001
R129 M42:BULK M27:BULK 0.001
R130 M42:BULK M30:BULK 0.001
R131 M42:BULK M29:BULK 0.001
R132 M42:BULK M32:BULK 0.001
R133 M42:BULK M31:BULK 0.001
R134 M42:BULK M36:BULK 0.001
R135 M42:BULK M35:BULK 0.001
R136 M42:BULK M34:BULK 0.001
R137 M42:BULK M33:BULK 0.001
R138 M42:BULK M40:BULK 0.001
R139 M42:BULK M39:BULK 0.001
R140 M42:BULK M38:BULK 0.001
R141 M42:BULK M37:BULK 0.001
R142 VDD M41:SRC 3.75474
R143 M30:SRC M41:SRC 6.80162e-10
R144 M30:SRC M29:SRC 0.001
R145 M32:SRC M41:SRC 5e-10
R146 M32:SRC M37:DRN 342.257
R147 M31:SRC M36:SRC 0.001
R148 M31:SRC M41:SRC 7.37374e-10
R149 M35:DRN M34:SRC 0.001
R150 M35:DRN M41:SRC 6.36364e-10
R151 M33:SRC M40:SRC 0.001
R152 M33:SRC M41:SRC 1.01515e-09
R153 M39:DRN M38:SRC 0.001
R154 M39:DRN M41:SRC 6.16601e-10
R155 M37:DRN M41:SRC 28.0442
R156 M41:SRC M42:DRN 0.001
R157 M26:DRN M23:SRC 6e-10
R158 N_16:1 N_16:3 20.1186
R159 N_16:1 M17:SRC 512.703
R160 N_16:1 M16:DRN 349.13
R161 N_16:1 M10:GATE 46.0358
R162 N_16:1 M9:GATE 137.142
R163 N_16:1 N_16:2 31.4452
R164 N_16:1 M40:GATE 66.96
R165 N_16:1 M39:GATE 163.515
R166 N_16:2 M9:GATE 135.203
R167 N_16:2 M8:GATE 56.16
R168 N_16:2 M7:GATE 83.6558
R169 N_16:2 M39:GATE 161.204
R170 N_16:2 M38:GATE 66.96
R171 N_16:2 M37:GATE 99.7434
R172 N_16:3 M17:SRC 20.0936
R173 N_16:3 M30:DRN 18
R174 N_16:3 M16:DRN 20.8168
R175 N_16:3 M29:DRN 18.4128
R176 M39:GATE M9:GATE 703.056
R177 M37:GATE M7:GATE 374.592
R178 M30:DRN M27:SRC 0.001
R179 M16:DRN M17:SRC 530.498
R180 M19:DRN M17:SRC 6.74817e-10
R181 N_8:1 N_8:5 15.1222
R182 N_8:1 M6:GATE 46.4965
R183 N_8:1 M5:GATE 139.717
R184 N_8:1 N_8:3 32.0357
R185 N_8:1 M36:GATE 66.96
R186 N_8:1 M35:GATE 166.586
R187 N_8:2 M17:GATE 45.84
R188 N_8:2 N_8:4 16.5733
R189 N_8:2 M1:DRN 1351.99
R190 N_8:2 N_8:5 42.1129
R191 N_8:2 M30:GATE 78.84
R192 N_8:3 M5:GATE 133.497
R193 N_8:3 M4:GATE 56.16
R194 N_8:3 M3:GATE 83.6558
R195 N_8:3 M35:GATE 159.169
R196 N_8:3 M34:GATE 66.96
R197 N_8:3 M33:GATE 99.7434
R198 N_8:4 M29:GATE 78.84
R199 N_8:4 M16:GATE 45.84
R200 N_8:4 M1:DRN 1272.46
R201 N_8:4 N_8:5 39.6356
R202 N_8:5 M32:DRN 9.56088
R203 N_8:5 M1:DRN 19.0848
R204 M35:GATE M5:GATE 694.183
R205 M33:GATE M3:GATE 374.592
R206 M32:DRN M31:DRN 0.001
R207 M1:DRN M2:DRN 0.001
R208 N_24:1 M19:SRC 157.609
R209 N_24:1 M28:SRC 75.6123
R210 N_24:1 N_24:2 17.3518
R211 N_24:1 M1:GATE 56.16
R212 N_24:1 M31:GATE 66.96
R213 N_24:2 M19:SRC 176.151
R214 N_24:2 M2:GATE 56.16
R215 N_24:2 M28:SRC 84.5079
R216 N_24:2 M32:GATE 66.96
R217 M28:SRC M19:SRC 35.5751
R218 M28:SRC M27:DRN 8.33333e-10
R219 M12:SRC M19:SRC 0.001
c_1 M13:SRC 0 1.79324e-19 
c_2 M23:DRN M14:DRN 9.56797e-19 
c_3 M23:DRN 0 1.35625e-19 
c_4 M26:GATE M14:DRN 3.08613e-18 
c_5 M26:GATE 0 9.90927e-19 
c_6 M24:DRN M23:DRN 1.85117e-18 
c_7 M24:DRN 0 9.72829e-19 
c_8 M15:GATE 0 1.58549e-20 
c_9 M13:DRN 0 2.09862e-17 
c_10 M24:GATE M13:DRN 5.03267e-18 
c_11 M24:GATE M26:GATE 4.14506e-20 
c_12 M24:GATE M24:DRN 2.80896e-17 
c_13 M24:GATE 0 3.73908e-18 
c_14 D M13:SRC 7.52876e-19 
c_15 D M13:DRN 1.94156e-18 
c_16 D M26:GATE 1.67194e-20 
c_17 D M24:DRN 1.17158e-16 
c_18 D 0 5.84871e-18 
c_19 M13:GATE M13:DRN 1.51097e-17 
c_20 M13:GATE M15:GATE 9.88517e-20 
c_21 M13:GATE M26:GATE 3.98761e-18 
c_22 M13:GATE 0 3.14613e-18 
c_23 M25:DRN D 6.00648e-18 
c_24 M25:DRN M13:SRC 2.32052e-18 
c_25 M25:DRN 0 8.18766e-20 
c_26 M41:GATE 0 1.92256e-17 
c_27 CP 0 1.17606e-18 
c_28 M20:GATE 0 7.80711e-18 
c_29 M28:DRN M13:DRN 1.7715e-16 
c_30 M28:DRN M23:DRN 2.17028e-20 
c_31 M28:DRN M26:GATE 2.92747e-17 
c_32 M28:DRN M24:DRN 5.2198e-21 
c_33 M28:DRN 0 3.9745e-20 
c_34 M15:DRN M13:DRN 2.81029e-17 
c_35 M15:DRN M23:DRN 2.07387e-18 
c_36 M15:DRN M15:GATE 1.12463e-17 
c_37 M15:DRN M26:GATE 8.86049e-18 
c_38 M15:DRN 0 6.11562e-18 
c_39 M12:DRN M13:DRN 1.06081e-20 
c_40 M12:DRN M15:GATE 1.02548e-17 
c_41 M12:DRN M24:DRN 4.73158e-18 
c_42 M12:DRN 0 3.10711e-20 
c_43 M23:GATE M26:GATE 3.19802e-18 
c_44 M23:GATE M24:DRN 1.97679e-17 
c_45 M23:GATE 0 7.60559e-18 
c_46 M14:GATE M13:DRN 9.46497e-19 
c_47 M14:GATE M15:GATE 2.03834e-19 
c_48 M14:GATE M24:DRN 2.25794e-17 
c_49 M14:GATE 0 1.0523e-17 
c_50 Q 0 2.77013e-17 
c_51 M36:DRN 0 7.58319e-18 
c_52 M34:DRN 0 5.55576e-18 
c_53 M3:DRN 0 8.45291e-19 
c_54 M5:SRC 0 1.25291e-18 
c_55 QN 0 3.09394e-17 
c_56 M40:DRN 0 6.13549e-18 
c_57 M38:DRN 0 1.137e-20 
c_58 M10:DRN 0 3.97013e-18 
c_59 M8:DRN 0 1.25964e-18 
c_60 M21:BULK M13:GATE 3.78331e-18 
c_61 M21:BULK M14:GATE 3.19753e-18 
c_62 M21:BULK M15:GATE 1.14928e-17 
c_63 M21:BULK M15:DRN 6.24908e-18 
c_64 M21:BULK D 7.55068e-18 
c_65 M21:BULK M20:GATE 1.14332e-17 
c_66 M21:BULK CP 2.29985e-18 
c_67 M21:BULK QN 3.48986e-18 
c_68 M9:DRN QN 7.80063e-18 
c_69 M9:DRN 0 2.37309e-18 
c_70 M3:SRC QN 6.90035e-20 
c_71 M3:SRC Q 6.90035e-20 
c_72 M3:SRC 0 3.49353e-18 
c_73 M5:DRN Q 2.74535e-18 
c_74 M5:DRN 0 2.37309e-18 
c_75 M1:SRC 0 3.32675e-18 
c_76 GND:1 M13:SRC 3.63255e-19 
c_77 GND:1 M13:GATE 5.07866e-18 
c_78 GND:1 M13:DRN 3.89032e-19 
c_79 GND:1 M14:GATE 5.42814e-19 
c_80 GND:1 M15:GATE 2.45275e-18 
c_81 GND:1 M15:DRN 5.63537e-18 
c_82 GND:1 M26:GATE 1.4915e-19 
c_83 GND:1 D 6.9574e-19 
c_84 GND:1 M20:GATE 6.64737e-18 
c_85 GND:1 CP 2.92763e-18 
c_86 GND:1 M5:SRC 1.31321e-18 
c_87 GND:1 Q 4.51158e-18 
c_88 GND:1 M3:DRN 1.13202e-18 
c_89 GND:1 M10:DRN 2.42006e-18 
c_90 GND:1 QN 1.27584e-16 
c_91 GND:1 M8:DRN 2.93241e-18 
c_92 GND:1 0 2.88775e-16 
c_93 GND CP 3.44941e-19 
c_94 GND 0 6.34448e-17 
c_95 M16:SRC 0 1.32823e-18 
c_96 M2:SRC 0 4.99629e-18 
c_97 M7:DRN M8:DRN 2.88574e-18 
c_98 M7:DRN QN 8.07835e-20 
c_99 M7:DRN 0 4.57628e-18 
c_100 M20:SRC M14:DRN 9.28648e-19 
c_101 M20:SRC M13:SRC 7.02121e-18 
c_102 M20:SRC M13:GATE 9.44091e-18 
c_103 M20:SRC M13:DRN 6.90899e-18 
c_104 M20:SRC M14:GATE 8.17413e-20 
c_105 M20:SRC M15:GATE 4.32215e-18 
c_106 M20:SRC M15:DRN 2.03772e-18 
c_107 M20:SRC M12:DRN 8.60658e-18 
c_108 M20:SRC M24:DRN 4.74451e-20 
c_109 M20:SRC D 2.53387e-19 
c_110 M20:SRC M28:DRN 9.02166e-20 
c_111 M20:SRC M20:GATE 2.02788e-17 
c_112 M20:SRC CP 2.36925e-19 
c_113 M20:SRC M36:DRN 4.42193e-20 
c_114 M20:SRC M5:SRC 8.80476e-18 
c_115 M20:SRC Q 1.93674e-18 
c_116 M20:SRC M34:DRN 4.42193e-20 
c_117 M20:SRC M3:DRN 8.80476e-18 
c_118 M20:SRC M10:DRN 1.13251e-17 
c_119 M20:SRC M40:DRN 4.42193e-20 
c_120 M20:SRC QN 2.63416e-18 
c_121 M20:SRC M8:DRN 1.13251e-17 
c_122 M20:SRC M38:DRN 4.42193e-20 
c_123 M20:SRC 0 1.44918e-16 
c_124 M18:SRC M13:GATE 1.84084e-18 
c_125 M18:SRC M13:DRN 3.44809e-19 
c_126 M18:SRC 0 1.41386e-18 
c_127 M14:SRC M15:DRN 5.21552e-18 
c_128 M14:SRC M13:DRN 1.44685e-20 
c_129 M14:SRC 0 8.24106e-20 
c_130 M15:SRC M13:SRC 1.64496e-20 
c_131 M15:SRC M13:GATE 1.91103e-18 
c_132 M15:SRC M13:DRN 5.90913e-18 
c_133 M15:SRC M14:GATE 1.85399e-17 
c_134 M15:SRC M23:GATE 1.42173e-21 
c_135 M15:SRC M15:GATE 1.36175e-17 
c_136 M15:SRC M15:DRN 4.39755e-18 
c_137 M15:SRC M26:GATE 8.4971e-20 
c_138 M15:SRC M12:DRN 6.26544e-18 
c_139 M15:SRC 0 6.14342e-18 
c_140 N_28:1 GND:1 3.08831e-17 
c_141 N_28:1 M20:SRC 7.21695e-18 
c_142 N_28:1 M15:GATE 6.23495e-19 
c_143 N_28:1 M15:DRN 1.73131e-20 
c_144 N_28:1 M18:SRC 1.10803e-17 
c_145 N_28:1 D 1.1357e-18 
c_146 N_28:1 M20:GATE 1.65581e-17 
c_147 N_28:1 M21:BULK 1.56315e-17 
c_148 N_28:1 CP 1.43755e-16 
c_149 N_28:1 M41:GATE 1.18662e-17 
c_150 N_28:1 0 1.13921e-18 
c_151 M22:GATE M14:DRN 1.05318e-18 
c_152 M22:GATE M20:SRC 4.59299e-21 
c_153 M22:GATE M23:GATE 1.04876e-17 
c_154 M22:GATE M15:DRN 1.48801e-18 
c_155 M22:GATE M26:GATE 3.26411e-18 
c_156 M22:GATE M24:GATE 4.15375e-18 
c_157 M22:GATE M24:DRN 2.28064e-17 
c_158 M22:GATE D 2.02136e-18 
c_159 M22:GATE M41:GATE 5.63658e-21 
c_160 M22:GATE 0 4.39569e-19 
c_161 M42:GATE M26:GATE 5.76831e-18 
c_162 M42:GATE M24:GATE 1.1305e-19 
c_163 M42:GATE M28:DRN 1.18449e-17 
c_164 M42:GATE M41:GATE 1.82088e-17 
c_165 M42:GATE 0 6.9543e-18 
c_166 M28:GATE M15:SRC 6.12787e-20 
c_167 M28:GATE M20:SRC 1.84098e-18 
c_168 M28:GATE M13:DRN 7.98827e-18 
c_169 M28:GATE M23:DRN 3.50791e-18 
c_170 M28:GATE M23:GATE 1.11272e-17 
c_171 M28:GATE M15:DRN 1.43165e-17 
c_172 M28:GATE M26:GATE 6.09624e-18 
c_173 M28:GATE M12:DRN 1.08291e-20 
c_174 M28:GATE M24:GATE 1.16426e-17 
c_175 M28:GATE M24:DRN 1.93924e-17 
c_176 M28:GATE D 5.56056e-19 
c_177 M28:GATE M28:DRN 1.84897e-17 
c_178 M28:GATE M25:DRN 5.06282e-18 
c_179 M28:GATE M21:BULK 4.27604e-18 
c_180 M28:GATE M41:GATE 2.24796e-18 
c_181 M28:GATE 0 9.76976e-18 
c_182 M19:GATE GND:1 8.01915e-19 
c_183 M19:GATE M20:SRC 1.87707e-18 
c_184 M19:GATE M14:GATE 1.23813e-20 
c_185 M19:GATE M15:GATE 1.24349e-21 
c_186 M19:GATE M15:DRN 3.9814e-21 
c_187 M19:GATE 0 3.40135e-17 
c_188 M41:DRN M41:GATE 1.68758e-17 
c_189 M41:DRN CP 1.70487e-17 
c_190 M41:DRN M20:SRC 6.43947e-20 
c_191 M41:DRN 0 4.98609e-18 
c_192 M21:GATE GND:1 4.92507e-18 
c_193 M21:GATE M20:SRC 1.4705e-17 
c_194 M21:GATE M13:SRC 1.8989e-18 
c_195 M21:GATE M13:GATE 1.84949e-19 
c_196 M21:GATE M18:SRC 4.34034e-18 
c_197 M21:GATE D 6.13612e-18 
c_198 M21:GATE M20:GATE 4.73132e-18 
c_199 M21:GATE 0 5.22746e-18 
c_200 M18:GATE M15:SRC 5.99972e-19 
c_201 M18:GATE GND:1 2.7053e-18 
c_202 M18:GATE M20:SRC 9.44106e-18 
c_203 M18:GATE M13:SRC 1.04059e-19 
c_204 M18:GATE M13:GATE 6.10479e-18 
c_205 M18:GATE M13:DRN 1.36697e-19 
c_206 M18:GATE M15:GATE 3.13176e-22 
c_207 M18:GATE M26:GATE 8.91908e-20 
c_208 M18:GATE M18:SRC 1.62166e-17 
c_209 M18:GATE M24:GATE 1.22711e-17 
c_210 M18:GATE D 2.07249e-19 
c_211 M18:GATE M20:GATE 1.94889e-19 
c_212 M18:GATE M21:BULK 9.26563e-19 
c_213 M18:GATE 0 2.34018e-17 
c_214 M20:DRN M20:SRC 8.37217e-18 
c_215 M20:DRN CP 3.06477e-17 
c_216 M20:DRN GND 1.37808e-20 
c_217 M20:DRN GND:1 1.21111e-18 
c_218 M20:DRN 0 1.72013e-18 
c_219 N_26:1 M14:DRN 4.37929e-18 
c_220 N_26:1 M15:SRC 1.05182e-17 
c_221 N_26:1 GND:1 2.52761e-16 
c_222 N_26:1 M20:SRC 6.23025e-17 
c_223 N_26:1 M18:GATE 5.78394e-18 
c_224 N_26:1 M13:SRC 3.74988e-18 
c_225 N_26:1 M13:GATE 9.73396e-19 
c_226 N_26:1 M13:DRN 2.44086e-17 
c_227 N_26:1 M14:GATE 1.29053e-17 
c_228 N_26:1 M14:SRC 1.53607e-19 
c_229 N_26:1 M23:GATE 4.22344e-17 
c_230 N_26:1 M15:GATE 3.48257e-17 
c_231 N_26:1 M26:GATE 2.50813e-17 
c_232 N_26:1 M12:DRN 2.36904e-18 
c_233 N_26:1 M28:GATE 8.86954e-19 
c_234 N_26:1 M18:SRC 1.46003e-18 
c_235 N_26:1 M24:GATE 1.84887e-18 
c_236 N_26:1 D 6.80731e-17 
c_237 N_26:1 M28:DRN 1.57326e-19 
c_238 N_26:1 M21:GATE 2.05529e-17 
c_239 N_26:1 M25:DRN 2.82308e-19 
c_240 N_26:1 N_28:1 1.38256e-16 
c_241 N_26:1 M21:BULK 2.87068e-17 
c_242 N_26:1 M19:GATE 2.61146e-17 
c_243 N_26:1 GND 4.45476e-19 
c_244 N_26:1 M42:GATE 3.16729e-17 
c_245 N_26:1 M22:GATE 2.83067e-19 
c_246 N_26:1 0 1.73854e-17 
c_247 M27:GATE M20:SRC 1.23468e-21 
c_248 M27:GATE M26:GATE 1.49665e-19 
c_249 M27:GATE M28:GATE 1.92679e-18 
c_250 M27:GATE M28:DRN 1.14154e-21 
c_251 M27:GATE 0 7.49065e-18 
c_252 M42:SRC M20:SRC 1.69111e-20 
c_253 M42:SRC M15:GATE 1.31735e-19 
c_254 M42:SRC M15:DRN 5.49695e-17 
c_255 M42:SRC M28:GATE 1.26511e-17 
c_256 M42:SRC M24:GATE 3.82504e-20 
c_257 M42:SRC M24:DRN 2.58685e-21 
c_258 M42:SRC D 1.17788e-20 
c_259 M42:SRC M28:DRN 3.24595e-22 
c_260 M42:SRC M25:DRN 6.25022e-19 
c_261 M42:SRC N_28:1 1.74505e-17 
c_262 M42:SRC M42:GATE 2.44428e-17 
c_263 M42:SRC M41:DRN 1.42676e-18 
c_264 M42:SRC M22:GATE 1.20974e-17 
c_265 M42:SRC 0 3.23742e-18 
c_266 M25:GATE M13:SRC 2.23749e-18 
c_267 M25:GATE M26:GATE 9.29895e-19 
c_268 M25:GATE M28:GATE 4.72059e-18 
c_269 M25:GATE M24:GATE 1.8472e-17 
c_270 M25:GATE M24:DRN 5.32531e-19 
c_271 M25:GATE D 2.439e-18 
c_272 M25:GATE M25:DRN 1.65973e-18 
c_273 M25:GATE M42:GATE 5.3475e-19 
c_274 M25:GATE M22:GATE 2.20203e-19 
c_275 M25:GATE 0 1.0397e-17 
c_276 M12:GATE M15:SRC 1.16188e-18 
c_277 M12:GATE GND:1 1.61263e-19 
c_278 M12:GATE M20:SRC 3.43448e-17 
c_279 M12:GATE M13:GATE 2.56878e-22 
c_280 M12:GATE M14:GATE 1.9015e-19 
c_281 M12:GATE M23:GATE 9.64936e-20 
c_282 M12:GATE M15:GATE 8.71728e-18 
c_283 M12:GATE M15:DRN 2.7938e-17 
c_284 M12:GATE M28:GATE 1.79685e-18 
c_285 M12:GATE M24:DRN 2.82007e-18 
c_286 M12:GATE M28:DRN 3.84668e-18 
c_287 M12:GATE M21:BULK 4.2553e-18 
c_288 M12:GATE M19:GATE 3.9596e-18 
c_289 M12:GATE 0 1.21496e-17 
c_290 M11:GATE M15:SRC 1.83147e-18 
c_291 M11:GATE GND:1 8.98152e-19 
c_292 M11:GATE M20:SRC 5.9556e-18 
c_293 M11:GATE M18:GATE 1.29245e-19 
c_294 M11:GATE M13:GATE 7.94137e-18 
c_295 M11:GATE M13:DRN 1.64306e-17 
c_296 M11:GATE M14:GATE 6.87194e-18 
c_297 M11:GATE M15:GATE 4.97014e-19 
c_298 M11:GATE M15:DRN 8.14433e-18 
c_299 M11:GATE M28:GATE 1.26883e-20 
c_300 M11:GATE M24:DRN 1.13578e-17 
c_301 M11:GATE D 3.64504e-18 
c_302 M11:GATE N_28:1 1.10485e-19 
c_303 M11:GATE M21:BULK 5.03908e-18 
c_304 M11:GATE M22:GATE 1.07112e-18 
c_305 M11:GATE 0 7.36541e-18 
c_306 M21:SRC GND:1 2.50811e-18 
c_307 M21:SRC M20:SRC 1.10546e-17 
c_308 M21:SRC M13:SRC 9.66101e-19 
c_309 M21:SRC M13:DRN 3.36393e-21 
c_310 M21:SRC M26:GATE 3.95212e-17 
c_311 M21:SRC M28:GATE 2.23264e-18 
c_312 M21:SRC M18:SRC 2.64708e-17 
c_313 M21:SRC D 4.53586e-20 
c_314 M21:SRC M20:DRN 9.42378e-19 
c_315 M21:SRC M21:GATE 7.98106e-18 
c_316 M21:SRC N_28:1 4.82373e-17 
c_317 M21:SRC M19:GATE 1.46055e-19 
c_318 M21:SRC 0 1.12455e-17 
c_319 VDD:1 M23:GATE 5.39271e-18 
c_320 VDD:1 M15:GATE 3.1959e-19 
c_321 VDD:1 M15:DRN 2.94703e-17 
c_322 VDD:1 M26:GATE 6.51529e-18 
c_323 VDD:1 M28:GATE 1.94613e-18 
c_324 VDD:1 N_26:1 3.05319e-19 
c_325 VDD:1 M24:GATE 1.28183e-18 
c_326 VDD:1 M24:DRN 5.59155e-17 
c_327 VDD:1 D 6.54089e-20 
c_328 VDD:1 M28:DRN 1.70915e-19 
c_329 VDD:1 M25:GATE 4.67406e-18 
c_330 VDD:1 N_28:1 5.90603e-19 
c_331 VDD:1 M42:SRC 5.14708e-19 
c_332 VDD:1 M42:GATE 5.69695e-18 
c_333 VDD:1 M22:GATE 1.72794e-18 
c_334 VDD:1 M27:GATE 2.11016e-19 
c_335 VDD:1 M36:DRN 8.02204e-19 
c_336 VDD:1 Q 2.4009e-19 
c_337 VDD:1 M34:DRN 2.61161e-20 
c_338 VDD:1 M40:DRN 3.12305e-18 
c_339 VDD:1 QN 4.09786e-17 
c_340 VDD:1 M8:DRN 1.29566e-19 
c_341 VDD:1 M38:DRN 5.60879e-18 
c_342 VDD:1 M41:GATE 7.22757e-19 
c_343 VDD:1 0 4.99443e-17 
c_344 M42:BULK M23:GATE 4.57778e-18 
c_345 M42:BULK M15:GATE 1.66115e-17 
c_346 M42:BULK M15:DRN 7.51315e-18 
c_347 M42:BULK M26:GATE 2.5134e-18 
c_348 M42:BULK M28:GATE 3.64562e-17 
c_349 M42:BULK N_26:1 1.61105e-17 
c_350 M42:BULK M24:GATE 2.26272e-18 
c_351 M42:BULK M24:DRN 3.65572e-18 
c_352 M42:BULK D 8.44044e-18 
c_353 M42:BULK M28:DRN 3.60128e-19 
c_354 M42:BULK M25:GATE 2.81188e-18 
c_355 M42:BULK M20:GATE 1.40623e-18 
c_356 M42:BULK N_28:1 6.8295e-18 
c_357 M42:BULK CP 3.09361e-18 
c_358 M42:BULK M42:GATE 5.03877e-18 
c_359 M42:BULK M22:GATE 1.10467e-17 
c_360 M42:BULK M27:GATE 4.133e-18 
c_361 M42:BULK M36:DRN 2.05433e-18 
c_362 M42:BULK Q 7.96554e-18 
c_363 M42:BULK M34:DRN 4.10201e-18 
c_364 M42:BULK M40:DRN 3.49234e-18 
c_365 M42:BULK QN 1.11619e-17 
c_366 M42:BULK M38:DRN 3.85789e-18 
c_367 M42:BULK M41:GATE 6.45901e-18 
c_368 VDD M23:GATE 1.16821e-18 
c_369 VDD M15:GATE 2.73829e-17 
c_370 VDD M15:DRN 1.7206e-17 
c_371 VDD M26:GATE 1.23046e-18 
c_372 VDD M28:GATE 7.46657e-17 
c_373 VDD N_26:1 4.62155e-17 
c_374 VDD M24:GATE 1.65875e-18 
c_375 VDD M24:DRN 1.60858e-18 
c_376 VDD D 2.8437e-18 
c_377 VDD M28:DRN 1.7911e-18 
c_378 VDD M25:GATE 9.44885e-19 
c_379 VDD N_28:1 2.85942e-17 
c_380 VDD M42:SRC 1.02529e-18 
c_381 VDD CP 1.18549e-18 
c_382 VDD M42:GATE 2.6513e-18 
c_383 VDD M41:DRN 1.10679e-18 
c_384 VDD M22:GATE 5.11565e-18 
c_385 VDD M27:GATE 1.94647e-18 
c_386 VDD M36:DRN 2.81065e-18 
c_387 VDD Q 9.44826e-17 
c_388 VDD M34:DRN 2.81065e-18 
c_389 VDD M40:DRN 2.81065e-18 
c_390 VDD QN 8.74e-17 
c_391 VDD M38:DRN 2.80996e-18 
c_392 VDD M41:GATE 9.00454e-18 
c_393 VDD 0 2.19741e-16 
c_394 M30:SRC M28:GATE 6.68189e-19 
c_395 M30:SRC M42:SRC 1.2322e-23 
c_396 M30:SRC 0 1.53659e-18 
c_397 M32:SRC M28:GATE 4.76795e-20 
c_398 M32:SRC M24:DRN 2.08641e-20 
c_399 M32:SRC M28:DRN 3.48112e-22 
c_400 M32:SRC M25:DRN 3.81897e-23 
c_401 M32:SRC M22:GATE 2.62568e-20 
c_402 M32:SRC M41:GATE 1.59073e-22 
c_403 M32:SRC 0 1.10261e-17 
c_404 M31:SRC Q 9.0373e-21 
c_405 M31:SRC 0 3.32871e-18 
c_406 M35:DRN Q 1.16562e-17 
c_407 M35:DRN 0 2.56554e-18 
c_408 M33:SRC QN 2.26367e-19 
c_409 M33:SRC Q 2.26367e-19 
c_410 M33:SRC 0 3.8091e-18 
c_411 M39:DRN QN 1.03274e-17 
c_412 M39:DRN 0 2.56554e-18 
c_413 M37:DRN M38:DRN 2.70806e-18 
c_414 M37:DRN QN 7.93306e-19 
c_415 M37:DRN M8:DRN 8.04549e-20 
c_416 M37:DRN 0 1.10183e-17 
c_417 M41:SRC M13:DRN 8.95128e-20 
c_418 M41:SRC M23:DRN 9.50272e-19 
c_419 M41:SRC M23:GATE 1.29619e-18 
c_420 M41:SRC M15:GATE 2.32487e-19 
c_421 M41:SRC M15:DRN 1.40253e-19 
c_422 M41:SRC M26:GATE 1.81361e-18 
c_423 M41:SRC M12:DRN 7.37055e-20 
c_424 M41:SRC M12:GATE 1.50365e-24 
c_425 M41:SRC M28:GATE 1.34401e-16 
c_426 M41:SRC M21:SRC 1.63435e-22 
c_427 M41:SRC M24:GATE 1.77533e-18 
c_428 M41:SRC M24:DRN 2.96264e-18 
c_429 M41:SRC D 3.38213e-20 
c_430 M41:SRC M28:DRN 5.82882e-18 
c_431 M41:SRC M20:DRN 5.33454e-20 
c_432 M41:SRC M25:GATE 1.71914e-18 
c_433 M41:SRC M25:DRN 2.74408e-18 
c_434 M41:SRC N_28:1 8.06989e-18 
c_435 M41:SRC M42:SRC 5.27484e-18 
c_436 M41:SRC CP 1.82928e-19 
c_437 M41:SRC M42:GATE 4.11521e-18 
c_438 M41:SRC M41:DRN 8.39526e-18 
c_439 M41:SRC M22:GATE 9.08623e-17 
c_440 M41:SRC M27:GATE 3.53576e-18 
c_441 M41:SRC M36:DRN 1.13591e-17 
c_442 M41:SRC M5:SRC 3.81007e-20 
c_443 M41:SRC Q 2.34025e-18 
c_444 M41:SRC M34:DRN 1.13591e-17 
c_445 M41:SRC M3:DRN 3.81007e-20 
c_446 M41:SRC M10:DRN 3.81007e-20 
c_447 M41:SRC M40:DRN 1.13591e-17 
c_448 M41:SRC QN 2.16968e-18 
c_449 M41:SRC M8:DRN 3.81007e-20 
c_450 M41:SRC M38:DRN 1.13591e-17 
c_451 M41:SRC M41:GATE 2.01808e-17 
c_452 M41:SRC 0 2.1369e-16 
c_453 M25:SRC M28:GATE 2.33535e-17 
c_454 M25:SRC N_26:1 2.19401e-18 
c_455 M25:SRC M24:GATE 2.54637e-18 
c_456 M25:SRC M24:DRN 2.00344e-19 
c_457 M25:SRC M28:DRN 1.36149e-19 
c_458 M25:SRC M21:GATE 2.82477e-18 
c_459 M25:SRC M25:GATE 2.33234e-17 
c_460 M25:SRC M42:SRC 3.14443e-17 
c_461 M25:SRC M42:GATE 1.30585e-18 
c_462 M25:SRC M22:GATE 2.4283e-18 
c_463 M25:SRC QN 4.02962e-19 
c_464 M25:SRC M41:GATE 1.99426e-19 
c_465 M25:SRC 0 1.95668e-18 
c_466 M26:DRN M13:DRN 1.30733e-17 
c_467 M26:DRN M23:GATE 2.11789e-17 
c_468 M26:DRN M15:DRN 6.59988e-19 
c_469 M26:DRN M26:GATE 1.1748e-17 
c_470 M26:DRN M12:DRN 8.32245e-19 
c_471 M26:DRN M28:GATE 1.31466e-20 
c_472 M26:DRN M24:DRN 2.34493e-18 
c_473 M26:DRN M28:DRN 9.95923e-19 
c_474 M26:DRN M25:DRN 7.30046e-21 
c_475 M26:DRN M42:GATE 8.36081e-18 
c_476 M26:DRN M22:GATE 1.7031e-18 
c_477 M26:DRN 0 3.93715e-18 
c_478 N_16:1 GND:1 1.14751e-18 
c_479 N_16:1 M20:SRC 3.66042e-19 
c_480 N_16:1 M41:SRC 4.01696e-19 
c_481 N_16:1 M42:BULK 8.10001e-19 
c_482 N_16:1 N_26:1 3.58037e-17 
c_483 N_16:1 M21:BULK 8.42778e-18 
c_484 N_16:1 Q 1.20505e-18 
c_485 N_16:1 M3:DRN 1.73716e-19 
c_486 N_16:1 M10:DRN 4.15512e-17 
c_487 N_16:1 M40:DRN 1.49115e-17 
c_488 N_16:1 M9:DRN 1.01575e-17 
c_489 N_16:1 M39:DRN 1.02252e-17 
c_490 N_16:1 QN 8.79101e-17 
c_491 N_16:1 M8:DRN 1.52448e-17 
c_492 N_16:1 M38:DRN 1.47549e-17 
c_493 N_16:1 VDD 6.05007e-19 
c_494 N_16:2 GND:1 7.41087e-18 
c_495 N_16:2 M20:SRC 1.63248e-19 
c_496 N_16:2 M42:BULK 2.86493e-18 
c_497 N_16:2 M21:BULK 8.11554e-18 
c_498 N_16:2 M10:DRN 9.95772e-18 
c_499 N_16:2 QN 3.15767e-17 
c_500 N_16:2 M8:DRN 2.95176e-17 
c_501 N_16:3 GND:1 2.18815e-16 
c_502 N_16:3 M20:SRC 6.20705e-17 
c_503 N_16:3 M41:SRC 3.48757e-18 
c_504 N_16:3 M42:BULK 5.11218e-18 
c_505 N_16:3 VDD:1 5.27887e-19 
c_506 N_16:3 N_26:1 1.60141e-17 
c_507 N_16:3 M21:BULK 1.31065e-17 
c_508 N_16:3 M27:GATE 9.47071e-18 
c_509 N_16:3 M30:SRC 3.14498e-18 
c_510 N_16:3 M16:SRC 3.01848e-18 
c_511 N_16:3 M2:SRC 2.5793e-18 
c_512 N_16:3 M1:SRC 3.20661e-18 
c_513 N_16:3 M5:SRC 5.42608e-18 
c_514 N_16:3 M5:DRN 2.11637e-18 
c_515 N_16:3 Q 1.26442e-16 
c_516 N_16:3 M3:DRN 5.76445e-18 
c_517 N_16:3 M3:SRC 6.68345e-18 
c_518 N_16:3 M33:SRC 3.2417e-18 
c_519 N_16:3 M10:DRN 2.29361e-18 
c_520 N_16:3 M40:DRN 1.19058e-18 
c_521 N_16:3 QN 7.43128e-17 
c_522 N_16:3 VDD 8.80588e-18 
c_523 N_16:3 0 7.53175e-18 
c_524 M40:GATE M41:SRC 9.0614e-18 
c_525 M40:GATE M42:BULK 3.22857e-18 
c_526 M40:GATE VDD:1 6.79106e-19 
c_527 M40:GATE Q 3.32213e-18 
c_528 M40:GATE M34:DRN 2.95269e-19 
c_529 M40:GATE M33:SRC 1.00916e-17 
c_530 M40:GATE M40:DRN 3.38972e-17 
c_531 M40:GATE M39:DRN 8.3293e-19 
c_532 M40:GATE QN 9.68949e-18 
c_533 M40:GATE VDD 7.62353e-18 
c_534 M40:GATE 0 8.97927e-19 
c_535 M39:GATE M41:SRC 9.49913e-18 
c_536 M39:GATE M42:BULK 3.77071e-19 
c_537 M39:GATE VDD:1 5.87395e-19 
c_538 M39:GATE Q 4.29482e-21 
c_539 M39:GATE M33:SRC 8.3293e-19 
c_540 M39:GATE M40:DRN 3.32546e-17 
c_541 M39:GATE M39:DRN 1.00916e-17 
c_542 M39:GATE QN 1.97601e-17 
c_543 M39:GATE M38:DRN 2.95269e-19 
c_544 M39:GATE VDD 7.35797e-18 
c_545 M38:GATE M41:SRC 9.49913e-18 
c_546 M38:GATE M42:BULK 5.0857e-18 
c_547 M38:GATE VDD:1 1.16292e-18 
c_548 M38:GATE M40:DRN 2.95269e-19 
c_549 M38:GATE M39:DRN 1.002e-17 
c_550 M38:GATE QN 2.04606e-17 
c_551 M38:GATE M38:DRN 3.34413e-17 
c_552 M38:GATE M37:DRN 3.2182e-20 
c_553 M38:GATE VDD 7.43949e-18 
c_554 M38:GATE 0 7.11157e-19 
c_555 M37:GATE M41:SRC 9.49797e-18 
c_556 M37:GATE M42:BULK 8.89374e-18 
c_557 M37:GATE VDD:1 6.73559e-18 
c_558 M37:GATE M39:DRN 1.12569e-18 
c_559 M37:GATE QN 1.13145e-17 
c_560 M37:GATE M8:DRN 7.07981e-18 
c_561 M37:GATE M38:DRN 3.279e-17 
c_562 M37:GATE M37:DRN 3.44923e-17 
c_563 M37:GATE VDD 7.93153e-18 
c_564 M37:GATE M7:DRN 1.59984e-18 
c_565 M37:GATE 0 5.51341e-19 
c_566 M30:DRN M20:SRC 2.87439e-22 
c_567 M30:DRN M41:SRC 8.79863e-18 
c_568 M30:DRN M42:BULK 2.101e-18 
c_569 M30:DRN N_26:1 7.41593e-19 
c_570 M30:DRN M42:SRC 6.99099e-23 
c_571 M30:DRN M25:SRC 2.91874e-20 
c_572 M30:DRN M27:GATE 2.32311e-17 
c_573 M30:DRN VDD 1.50711e-18 
c_574 M30:DRN 0 7.13267e-19 
c_575 M29:DRN M20:SRC 5.35969e-20 
c_576 M29:DRN M41:SRC 7.97399e-18 
c_577 M29:DRN VDD:1 1.81287e-19 
c_578 M29:DRN M32:SRC 2.97237e-17 
c_579 M29:DRN VDD 1.24192e-18 
c_580 M29:DRN 0 4.25769e-18 
c_581 M8:GATE M21:BULK 4.37806e-18 
c_582 M8:GATE QN 2.24691e-19 
c_583 M8:GATE GND:1 4.68162e-18 
c_584 M8:GATE M8:DRN 2.07716e-17 
c_585 M8:GATE M7:DRN 4.16913e-20 
c_586 M8:GATE M20:SRC 1.94243e-17 
c_587 M10:GATE M21:BULK 1.73848e-18 
c_588 M10:GATE QN 2.88218e-19 
c_589 M10:GATE GND:1 3.41962e-18 
c_590 M10:GATE M10:DRN 1.199e-17 
c_591 M10:GATE M20:SRC 2.05767e-17 
c_592 M10:GATE 0 3.26394e-18 
c_593 M9:GATE M21:BULK 5.67825e-18 
c_594 M9:GATE QN 3.43328e-18 
c_595 M9:GATE GND:1 3.1418e-18 
c_596 M9:GATE M10:DRN 1.921e-17 
c_597 M9:GATE M8:DRN 2.02241e-19 
c_598 M9:GATE M20:SRC 2.09991e-17 
c_599 M7:GATE M21:BULK 9.58451e-18 
c_600 M7:GATE GND:1 5.32245e-18 
c_601 M7:GATE M8:DRN 1.02359e-17 
c_602 M7:GATE M7:DRN 3.35994e-17 
c_603 M7:GATE M20:SRC 1.12087e-17 
c_604 M16:DRN GND:1 1.90239e-18 
c_605 M16:DRN M20:SRC 1.11767e-17 
c_606 M16:DRN M41:SRC 5.05586e-20 
c_607 M16:DRN N_26:1 3.76198e-17 
c_608 M16:DRN M2:SRC 2.22789e-17 
c_609 M16:DRN 0 8.74645e-18 
c_610 M19:DRN N_26:1 1.5188e-18 
c_611 M19:DRN GND:1 3.7667e-20 
c_612 M19:DRN M12:GATE 1.1639e-18 
c_613 M19:DRN M20:SRC 9.16706e-18 
c_614 M19:DRN 0 5.588e-18 
c_615 M17:SRC GND:1 1.14201e-18 
c_616 M17:SRC M20:SRC 1.77302e-18 
c_617 M17:SRC M41:SRC 2.91529e-22 
c_618 M17:SRC M12:GATE 2.29556e-21 
c_619 M17:SRC N_26:1 3.53517e-17 
c_620 M17:SRC 0 1.31842e-17 
c_621 N_8:1 GND:1 5.27473e-19 
c_622 N_8:1 M20:SRC 6.4801e-19 
c_623 N_8:1 M41:SRC 4.02451e-19 
c_624 N_8:1 M21:BULK 4.31172e-18 
c_625 N_8:1 N_16:3 2.19448e-17 
c_626 N_8:1 M36:DRN 1.50108e-17 
c_627 N_8:1 M5:SRC 2.64575e-17 
c_628 N_8:1 M5:DRN 1.01687e-17 
c_629 N_8:1 M35:DRN 1.02252e-17 
c_630 N_8:1 Q 4.06923e-17 
c_631 N_8:1 M34:DRN 1.49144e-17 
c_632 N_8:1 M3:DRN 1.63103e-17 
c_633 N_8:1 N_16:1 9.92522e-18 
c_634 N_8:1 VDD 6.05007e-19 
c_635 N_8:2 GND:1 9.98328e-19 
c_636 N_8:2 M20:SRC 5.86416e-19 
c_637 N_8:2 M41:SRC 4.6379e-19 
c_638 N_8:2 M42:BULK 3.57472e-18 
c_639 N_8:2 M21:BULK 7.15664e-18 
c_640 N_8:2 N_16:3 2.46993e-17 
c_641 N_8:2 M17:SRC 6.2888e-18 
c_642 N_8:2 M30:SRC 5.70555e-18 
c_643 N_8:2 M16:SRC 1.72072e-17 
c_644 N_8:2 0 2.44764e-17 
c_645 N_8:3 GND:1 1.58242e-18 
c_646 N_8:3 M20:SRC 1.48737e-19 
c_647 N_8:3 M42:BULK 9.27697e-19 
c_648 N_8:3 M21:BULK 6.95309e-18 
c_649 N_8:3 GND 7.16399e-19 
c_650 N_8:3 N_16:3 1.93461e-17 
c_651 N_8:3 M5:SRC 5.47033e-18 
c_652 N_8:3 Q 1.66044e-17 
c_653 N_8:3 M3:DRN 5.94184e-18 
c_654 N_8:3 N_16:1 3.45248e-18 
c_655 N_8:3 N_16:2 1.92173e-19 
c_656 N_8:3 M40:GATE 1.83676e-18 
c_657 N_8:4 M20:SRC 2.09883e-20 
c_658 N_8:4 M21:BULK 1.15878e-18 
c_659 N_8:4 N_16:3 8.03337e-18 
c_660 N_8:4 M17:SRC 1.274e-19 
c_661 N_8:4 M16:DRN 5.68652e-18 
c_662 N_8:4 M32:SRC 5.03408e-18 
c_663 N_8:4 M5:SRC 6.52692e-20 
c_664 N_8:4 Q 3.31894e-19 
c_665 N_8:4 0 3.33243e-18 
c_666 N_8:5 GND:1 4.4593e-18 
c_667 N_8:5 M20:SRC 4.21377e-18 
c_668 N_8:5 M41:SRC 1.23928e-18 
c_669 N_8:5 M42:BULK 1.01976e-17 
c_670 N_8:5 VDD:1 1.12026e-17 
c_671 N_8:5 GND 2.14692e-18 
c_672 N_8:5 N_16:3 2.09409e-16 
c_673 N_8:5 M30:DRN 8.44119e-20 
c_674 N_8:5 M16:DRN 2.99377e-18 
c_675 N_8:5 M29:DRN 1.89575e-18 
c_676 N_8:5 M2:SRC 5.49915e-18 
c_677 N_8:5 M32:SRC 1.32522e-18 
c_678 N_8:5 M1:SRC 4.34686e-18 
c_679 N_8:5 M31:SRC 5.75773e-18 
c_680 N_8:5 M36:DRN 1.4041e-18 
c_681 N_8:5 M5:SRC 1.41295e-18 
c_682 N_8:5 Q 1.02248e-16 
c_683 N_8:5 VDD 4.3609e-17 
c_684 N_8:5 0 4.00936e-18 
c_685 M36:GATE M41:SRC 9.49913e-18 
c_686 M36:GATE M42:BULK 3.78241e-18 
c_687 M36:GATE VDD:1 6.51229e-19 
c_688 M36:GATE M31:SRC 1.01282e-17 
c_689 M36:GATE M36:DRN 3.56194e-17 
c_690 M36:GATE M35:DRN 8.3293e-19 
c_691 M36:GATE Q 7.53553e-18 
c_692 M36:GATE VDD 6.93035e-18 
c_693 M36:GATE 0 5.25243e-19 
c_694 M35:GATE M41:SRC 9.49913e-18 
c_695 M35:GATE M42:BULK 5.23585e-18 
c_696 M35:GATE VDD:1 5.87395e-19 
c_697 M35:GATE M31:SRC 8.3293e-19 
c_698 M35:GATE M36:DRN 3.32286e-17 
c_699 M35:GATE M35:DRN 1.00916e-17 
c_700 M35:GATE Q 1.89391e-17 
c_701 M35:GATE M34:DRN 2.95269e-19 
c_702 M35:GATE VDD 7.35797e-18 
c_703 M34:GATE M41:SRC 9.49913e-18 
c_704 M34:GATE M42:BULK 5.47764e-18 
c_705 M34:GATE VDD:1 6.79106e-19 
c_706 M34:GATE M36:DRN 2.95269e-19 
c_707 M34:GATE M35:DRN 1.00916e-17 
c_708 M34:GATE Q 2.06776e-17 
c_709 M34:GATE M34:DRN 3.32605e-17 
c_710 M34:GATE M33:SRC 8.3293e-19 
c_711 M34:GATE VDD 7.33237e-18 
c_712 M34:GATE M40:GATE 3.98856e-19 
c_713 M34:GATE 0 5.95811e-19 
c_714 M33:GATE M41:SRC 9.0614e-18 
c_715 M33:GATE M42:BULK 4.02274e-18 
c_716 M33:GATE VDD:1 5.87395e-19 
c_717 M33:GATE N_16:3 1.28248e-18 
c_718 M33:GATE M35:DRN 8.3293e-19 
c_719 M33:GATE Q 1.18438e-17 
c_720 M33:GATE M34:DRN 3.38457e-17 
c_721 M33:GATE M33:SRC 1.00916e-17 
c_722 M33:GATE N_16:1 5.48084e-18 
c_723 M33:GATE N_16:2 3.30984e-20 
c_724 M33:GATE VDD 7.64913e-18 
c_725 M33:GATE M40:GATE 1.99018e-17 
c_726 M33:GATE M39:GATE 2.33063e-19 
c_727 M33:GATE 0 1.99992e-18 
c_728 M30:GATE M41:SRC 8.62966e-18 
c_729 M30:GATE M42:BULK 1.17995e-17 
c_730 M30:GATE VDD:1 1.3976e-18 
c_731 M30:GATE N_16:3 6.54049e-18 
c_732 M30:GATE M30:DRN 1.77285e-17 
c_733 M30:GATE M30:SRC 1.07628e-17 
c_734 M30:GATE M29:DRN 1.274e-19 
c_735 M30:GATE M32:SRC 1.04673e-18 
c_736 M30:GATE VDD 5.90571e-18 
c_737 M30:GATE 0 8.44549e-18 
c_738 M29:GATE M41:SRC 8.87307e-18 
c_739 M29:GATE M42:BULK 3.67505e-18 
c_740 M29:GATE VDD:1 1.11267e-18 
c_741 M29:GATE N_16:3 1.02937e-17 
c_742 M29:GATE M30:DRN 1.274e-19 
c_743 M29:GATE M30:SRC 5.26149e-18 
c_744 M29:GATE M29:DRN 1.66937e-17 
c_745 M29:GATE M32:SRC 3.9349e-18 
c_746 M29:GATE VDD 5.87661e-18 
c_747 M29:GATE 0 6.39373e-19 
c_748 M32:DRN M20:SRC 2.68579e-20 
c_749 M32:DRN M41:SRC 1.10518e-17 
c_750 M32:DRN M42:BULK 2.45436e-18 
c_751 M32:DRN VDD:1 3.35973e-20 
c_752 M32:DRN M30:SRC 2.07592e-22 
c_753 M32:DRN M29:DRN 7.1976e-20 
c_754 M32:DRN M36:DRN 5.78741e-20 
c_755 M32:DRN Q 3.42487e-19 
c_756 M32:DRN VDD 2.21153e-18 
c_757 M32:DRN 0 1.12877e-17 
c_758 M4:GATE N_16:1 2.64425e-19 
c_759 M4:GATE Q 1.31243e-19 
c_760 M4:GATE N_16:3 1.23056e-19 
c_761 M4:GATE M21:BULK 5.23502e-18 
c_762 M4:GATE M10:GATE 3.89664e-19 
c_763 M4:GATE GND:1 3.12894e-18 
c_764 M4:GATE M3:DRN 1.29107e-17 
c_765 M4:GATE M20:SRC 2.0999e-17 
c_766 M4:GATE 0 7.43145e-20 
c_767 M3:GATE GND:1 3.41962e-18 
c_768 M3:GATE M20:SRC 2.05767e-17 
c_769 M3:GATE M21:BULK 5.13787e-18 
c_770 M3:GATE N_16:3 1.69712e-19 
c_771 M3:GATE Q 6.56216e-20 
c_772 M3:GATE M3:DRN 1.56681e-17 
c_773 M3:GATE M10:GATE 4.53526e-18 
c_774 M3:GATE N_16:1 7.64371e-18 
c_775 M3:GATE M9:GATE 3.89664e-19 
c_776 M3:GATE 0 6.08516e-19 
c_777 M17:GATE N_16:3 7.73192e-19 
c_778 M17:GATE M21:BULK 3.77669e-18 
c_779 M17:GATE GND:1 2.12493e-18 
c_780 M17:GATE M16:DRN 1.274e-19 
c_781 M17:GATE M17:SRC 1.27172e-17 
c_782 M17:GATE M20:SRC 1.55612e-17 
c_783 M17:GATE 0 5.07973e-18 
c_784 M16:GATE N_16:3 1.54038e-18 
c_785 M16:GATE GND:1 2.0695e-18 
c_786 M16:GATE M16:DRN 1.1164e-17 
c_787 M16:GATE M2:SRC 3.08417e-18 
c_788 M16:GATE M20:SRC 1.28267e-17 
c_789 M16:GATE 0 1.01504e-18 
c_790 M6:GATE Q 5.90535e-19 
c_791 M6:GATE N_16:3 1.10903e-19 
c_792 M6:GATE M21:BULK 7.39364e-19 
c_793 M6:GATE GND:1 3.12894e-18 
c_794 M6:GATE M5:SRC 8.57032e-18 
c_795 M6:GATE M20:SRC 2.0999e-17 
c_796 M6:GATE 0 2.35313e-18 
c_797 M5:GATE GND:1 3.12894e-18 
c_798 M5:GATE M20:SRC 2.0999e-17 
c_799 M5:GATE M21:BULK 5.57264e-18 
c_800 M5:GATE N_16:3 1.23056e-19 
c_801 M5:GATE M5:SRC 1.05875e-17 
c_802 M5:GATE Q 4.19678e-18 
c_803 M5:GATE M3:DRN 1.64411e-19 
c_804 M1:DRN GND:1 1.4027e-18 
c_805 M1:DRN M20:SRC 8.6302e-18 
c_806 M1:DRN M41:SRC 1.93613e-20 
c_807 M1:DRN N_16:3 5.50253e-18 
c_808 M1:DRN M16:DRN 4.79976e-20 
c_809 M1:DRN M5:SRC 4.34055e-20 
c_810 M1:DRN Q 1.06087e-17 
c_811 M1:DRN 0 3.74783e-19 
c_812 N_24:1 GND:1 5.27473e-19 
c_813 N_24:1 M20:SRC 6.26687e-19 
c_814 N_24:1 M42:BULK 3.63294e-19 
c_815 N_24:1 N_26:1 2.52766e-17 
c_816 N_24:1 M29:GATE 3.69465e-20 
c_817 N_24:1 M21:BULK 2.44743e-18 
c_818 N_24:1 N_16:3 6.10989e-18 
c_819 N_24:1 N_8:2 8.21033e-21 
c_820 N_24:1 N_8:4 6.77706e-18 
c_821 N_24:1 M16:GATE 4.39542e-20 
c_822 N_24:1 M16:DRN 8.12425e-21 
c_823 N_24:1 M32:DRN 2.81582e-18 
c_824 N_24:1 M1:DRN 1.24606e-18 
c_825 N_24:1 N_8:5 8.20541e-17 
c_826 N_24:1 N_8:1 1.61969e-17 
c_827 N_24:1 N_8:3 3.69776e-19 
c_828 N_24:1 N_16:1 1.56818e-21 
c_829 N_24:1 M37:DRN 2.27259e-20 
c_830 N_24:1 M36:GATE 1.9401e-18 
c_831 N_24:1 M38:GATE 5.25367e-20 
c_832 N_24:1 M37:GATE 4.04e-20 
c_833 N_24:1 0 7.82522e-18 
c_834 N_24:2 M20:SRC 4.65049e-18 
c_835 N_24:2 M41:SRC 9.47259e-21 
c_836 N_24:2 M42:BULK 3.43823e-18 
c_837 N_24:2 M28:GATE 2.55329e-20 
c_838 N_24:2 M29:GATE 1.42334e-19 
c_839 N_24:2 M21:BULK 7.07079e-18 
c_840 N_24:2 N_16:3 6.80906e-18 
c_841 N_24:2 N_8:2 2.00232e-18 
c_842 N_24:2 M17:GATE 2.96212e-20 
c_843 N_24:2 N_8:4 1.12317e-18 
c_844 N_24:2 M16:GATE 6.25074e-19 
c_845 N_24:2 M16:DRN 1.02232e-18 
c_846 N_24:2 M32:DRN 1.45466e-17 
c_847 N_24:2 M1:DRN 1.66325e-17 
c_848 N_24:2 N_8:5 1.26231e-16 
c_849 N_24:2 N_8:1 1.11369e-17 
c_850 N_24:2 N_16:1 6.58635e-21 
c_851 N_24:2 M30:GATE 4.83816e-20 
c_852 N_24:2 0 2.17325e-18 
c_853 M32:GATE M41:SRC 9.06012e-18 
c_854 M32:GATE M42:BULK 4.89175e-18 
c_855 M32:GATE VDD:1 2.73307e-18 
c_856 M32:GATE M28:GATE 3.13636e-22 
c_857 M32:GATE M29:GATE 6.08943e-19 
c_858 M32:GATE N_16:3 1.45043e-18 
c_859 M32:GATE N_8:4 4.72943e-19 
c_860 M32:GATE M29:DRN 1.05797e-18 
c_861 M32:GATE M32:SRC 2.06798e-17 
c_862 M32:GATE M32:DRN 3.34968e-17 
c_863 M32:GATE M31:SRC 8.3293e-19 
c_864 M32:GATE N_8:5 5.96106e-18 
c_865 M32:GATE VDD 5.49396e-18 
c_866 M32:GATE M30:GATE 6.00296e-20 
c_867 M32:GATE M36:GATE 2.66618e-19 
c_868 M32:GATE 0 8.58923e-19 
c_869 M31:GATE M41:SRC 9.28177e-18 
c_870 M31:GATE M42:BULK 4.81096e-18 
c_871 M31:GATE VDD:1 9.32327e-19 
c_872 M31:GATE M29:GATE 4.45018e-20 
c_873 M31:GATE M29:DRN 4.51347e-22 
c_874 M31:GATE M32:SRC 1.47578e-18 
c_875 M31:GATE M32:DRN 3.57754e-17 
c_876 M31:GATE M31:SRC 1.00916e-17 
c_877 M31:GATE N_8:5 1.05207e-17 
c_878 M31:GATE VDD 5.63475e-18 
c_879 M31:GATE M36:GATE 1.91327e-17 
c_880 M31:GATE M35:GATE 2.33063e-19 
c_881 M31:GATE 0 1.3203e-18 
c_882 M28:SRC M20:SRC 1.08385e-19 
c_883 M28:SRC M41:SRC 5.93024e-17 
c_884 M28:SRC M42:BULK 1.19618e-17 
c_885 M28:SRC M14:GATE 5.13327e-17 
c_886 M28:SRC VDD:1 2.79871e-18 
c_887 M28:SRC M15:DRN 2.38122e-17 
c_888 M28:SRC M26:DRN 3.9065e-20 
c_889 M28:SRC M12:GATE 1.97201e-18 
c_890 M28:SRC M28:GATE 2.12604e-17 
c_891 M28:SRC N_26:1 3.4445e-17 
c_892 M28:SRC M29:GATE 9.90107e-18 
c_893 M28:SRC M28:DRN 4.4103e-17 
c_894 M28:SRC M21:BULK 3.83035e-18 
c_895 M28:SRC M19:GATE 4.92436e-17 
c_896 M28:SRC M25:SRC 3.77922e-20 
c_897 M28:SRC M27:GATE 4.89819e-17 
c_898 M28:SRC N_16:3 3.29326e-19 
c_899 M28:SRC N_8:2 1.41699e-18 
c_900 M28:SRC M30:DRN 1.30206e-17 
c_901 M28:SRC M30:SRC 2.37308e-18 
c_902 M28:SRC N_8:4 2.02132e-19 
c_903 M28:SRC M29:DRN 6.62437e-18 
c_904 M28:SRC M32:SRC 1.14647e-17 
c_905 M28:SRC M32:DRN 1.44397e-18 
c_906 M28:SRC VDD 1.24761e-16 
c_907 M28:SRC M30:GATE 9.07401e-18 
c_908 M28:SRC 0 3.77177e-18 
c_909 M1:GATE N_8:5 2.25248e-19 
c_910 M1:GATE N_16:3 1.12618e-19 
c_911 M1:GATE M21:BULK 3.57934e-18 
c_912 M1:GATE M6:GATE 4.30807e-18 
c_913 M1:GATE M5:GATE 2.84919e-19 
c_914 M1:GATE GND:1 3.27428e-18 
c_915 M1:GATE GND 6.82572e-19 
c_916 M1:GATE M1:DRN 1.77266e-17 
c_917 M1:GATE M20:SRC 2.07078e-17 
c_918 M2:GATE M15:SRC 3.18147e-22 
c_919 M2:GATE GND:1 3.13604e-18 
c_920 M2:GATE M20:SRC 2.77653e-17 
c_921 M2:GATE M12:GATE 5.87304e-20 
c_922 M2:GATE M21:BULK 1.16919e-18 
c_923 M2:GATE N_16:3 1.27419e-19 
c_924 M2:GATE M16:GATE 6.28642e-20 
c_925 M2:GATE M1:DRN 1.50959e-17 
c_926 M2:GATE N_8:5 1.65965e-19 
c_927 M2:GATE M6:GATE 2.12819e-19 
c_928 M2:GATE N_8:1 6.29771e-20 
c_929 M2:GATE 0 1.92129e-19 
c_930 M12:SRC M15:SRC 1.57973e-19 
c_931 M12:SRC M20:SRC 4.55846e-18 
c_932 M12:SRC M41:SRC 2.87819e-19 
c_933 M12:SRC M14:SRC 7.23426e-21 
c_934 M12:SRC M15:DRN 1.01629e-18 
c_935 M12:SRC M12:GATE 2.24361e-18 
c_936 M12:SRC M28:GATE 1.39655e-17 
c_937 M12:SRC N_26:1 2.25995e-17 
c_938 M12:SRC M28:DRN 1.63835e-18 
c_939 M12:SRC M19:GATE 1.44468e-18 
c_940 M12:SRC M27:GATE 1.06164e-19 
c_941 M12:SRC M19:DRN 1.15072e-18 
c_942 M12:SRC M17:GATE 7.05641e-19 
c_943 M12:SRC M16:SRC 1.49016e-20 
c_944 M12:SRC M2:SRC 3.41203e-22 
c_945 M19:SRC M15:SRC 3.098e-22 
c_946 M19:SRC M20:SRC 7.84968e-19 
c_947 M19:SRC M41:SRC 2.64601e-20 
c_948 M19:SRC M14:GATE 1.8584e-18 
c_949 M19:SRC M14:SRC 5.43879e-20 
c_950 M19:SRC M15:DRN 9.39719e-19 
c_951 M19:SRC M12:GATE 1.30027e-17 
c_952 M19:SRC N_26:1 7.98161e-17 
c_953 M19:SRC M28:DRN 2.28785e-21 
c_954 M19:SRC M19:GATE 1.59234e-17 
c_955 M19:SRC M19:DRN 1.19898e-18 
c_956 M19:SRC N_16:3 1.45821e-16 
c_957 M19:SRC M17:SRC 9.31833e-19 
c_958 M19:SRC N_8:2 3.2211e-20 
c_959 M19:SRC M16:SRC 7.50637e-21 
c_960 M19:SRC 0 2.84565e-20 

.ENDS
