
.subckt MUX4D1  I0 I1 I2 I3 S0 S1 Z
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.03483p as=0.03807p l=0.09u nrd=0.478 nrs=0.527 pd=0.5283u ps=0.5544u sa=1.449e-06 sb=2.835e-06 w=0.27u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.11664p as=0.10206p l=0.09u nrd=0.4 nrs=0.35 pd=1.512u ps=0.918u sa=2.16e-07 sb=1.4049e-06 w=0.54u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK nch ad=0.06885p as=0.11259p l=0.09u nrd=0.236 nrs=0.387 pd=0.8847u ps=1.3437u sa=5.85e-07 sb=3.312e-07 w=0.54u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.08424p as=0.04698p l=0.09u nrd=0.511 nrs=0.289 pd=1.224u ps=0.639u sa=2.07e-07 sb=5.58e-07 w=0.405u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.05427p as=0.081p l=0.09u nrd=0.74 nrs=1.111 pd=0.612u ps=0.756u sa=2.934e-06 sb=1.35e-06 w=0.27u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.12312p as=0.06966p l=0.09u nrd=0.421 nrs=0.239 pd=1.107u ps=1.0557u sa=2.826e-07 sb=1.1835e-06 w=0.54u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.05751p as=0.06642p l=0.09u nrd=0.351 nrs=0.403 pd=0.8316u ps=0.7173u sa=1.071e-06 sb=4.41e-07 w=0.405u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.10206p as=0.08829p l=0.09u nrd=0.35 nrs=0.302 pd=0.918u ps=0.9567u sa=6.84e-07 sb=6.597e-07 w=0.54u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK nch ad=0.0567p as=0.05832p l=0.09u nrd=0.774 nrs=0.8 pd=0.6723u ps=0.972u sa=4.068e-06 sb=2.16e-07 w=0.27u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.1134p as=0.04698p l=0.09u nrd=0.692 nrs=0.289 pd=1.476u ps=0.639u sa=5.31e-07 sb=2.34e-07 w=0.405u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.0972p as=0.11178p l=0.09u nrd=0.334 nrs=0.383 pd=1.764u ps=1.494u sa=1.44e-07 sb=2.07e-07 w=0.54u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.081p as=0.05184p l=0.09u nrd=0.493 nrs=0.314 pd=0.918u ps=0.6633u sa=7.722e-07 sb=7.443e-07 w=0.405u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.12312p as=0.162p l=0.09u nrd=0.421 nrs=0.556 pd=1.107u ps=1.512u sa=9.549e-07 sb=5.553e-07 w=0.54u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK pch ad=0.11178p as=0.13122p l=0.09u nrd=0.216 nrs=0.254 pd=1.2942u ps=1.224u sa=3.744e-07 sb=8.766e-07 w=0.72u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK pch ad=0.1053p as=0.05265p l=0.09u nrd=0.52 nrs=0.26 pd=1.368u ps=0.684u sa=2.79e-06 sb=2.34e-07 w=0.45u 
MM23 M23:DRN M23:GATE M23:SRC M23:BULK pch ad=0.17577p as=0.14904p l=0.09u nrd=0.339 nrs=0.287 pd=2.25u ps=1.854u sa=2.07e-07 sb=2.07e-07 w=0.72u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK pch ad=0.07776p as=0.0648p l=0.09u nrd=0.6 nrs=0.498 pd=1.152u ps=0.828u sa=5.4e-07 sb=2.16e-07 w=0.36u 
MM25 M25:DRN M25:GATE M25:SRC M25:BULK pch ad=0.11502p as=0.1215p l=0.09u nrd=0.222 nrs=0.235 pd=1.188u ps=1.3383u sa=5.76e-07 sb=3.897e-07 w=0.72u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK pch ad=0.08181p as=0.0729p l=0.09u nrd=0.438 nrs=0.391 pd=0.81u ps=0.8028u sa=1.017e-06 sb=2.151e-06 w=0.432u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK pch ad=0.06642p as=0.12636p l=0.09u nrd=0.228 nrs=0.433 pd=0.9018u ps=1.548u sa=3.447e-07 sb=2.34e-07 w=0.54u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK pch ad=0.13122p as=0.09315p l=0.09u nrd=0.254 nrs=0.18 pd=1.224u ps=1.1745u sa=1.0233e-06 sb=3.699e-07 w=0.72u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK pch ad=0.11583p as=0.06075p l=0.09u nrd=0.473 nrs=0.248 pd=1.458u ps=0.8262u sa=2.34e-07 sb=3.861e-07 w=0.495u 
MM24 M24:DRN M24:GATE M24:SRC M24:BULK pch ad=0.15552p as=0.11502p l=0.09u nrd=0.3 nrs=0.222 pd=1.872u ps=1.188u sa=2.16e-07 sb=1.0395e-06 w=0.72u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK pch ad=0.05265p as=0.05832p l=0.09u nrd=0.26 nrs=0.288 pd=0.684u ps=0.7335u sa=2.4426e-06 sb=5.58e-07 w=0.45u 
MM26 M26:DRN M26:GATE M26:SRC M26:BULK pch ad=0.16848p as=0.12879p l=0.09u nrd=0.325 nrs=0.249 pd=1.908u ps=1.656u sa=2.34e-07 sb=2.835e-07 w=0.72u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK pch ad=0.08181p as=0.06723p l=0.09u nrd=0.438 nrs=0.36 pd=0.81u ps=0.7767u sa=1.485e-06 sb=1.683e-06 w=0.432u 
R1 M25:SRC M11:SRC 36.3919
R2 M25:SRC M18:SRC 0.001
R3 M11:SRC M8:SRC 0.001
R4 M22:GATE I2 93.2367
R5 M22:GATE M7:GATE 305.443
R6 I2 M7:GATE 76.4373
R7 M21:GATE M6:GATE 342.936
R8 M21:GATE I0 89.7424
R9 I0 M6:GATE 86.8339
R10 M25:GATE I1 92.6419
R11 M25:GATE M11:GATE 299.553
R12 I1 M11:GATE 75.77
R13 M5:GATE S0 391.453
R14 M5:GATE M19:GATE 10896.8
R15 M5:GATE M17:GATE 816.426
R16 M24:GATE S0 93.2367
R17 M24:GATE M10:GATE 305.443
R18 M17:GATE S0 61.4137
R19 M17:GATE M19:GATE 1709.57
R20 M19:GATE S0 55.0208
R21 M19:GATE M8:GATE 141.36
R22 S0 M10:GATE 76.4373
R23 M21:DRN M6:SRC 36.436
R24 M21:DRN M19:SRC 0.001
R25 M6:SRC M9:DRN 0.001
R26 M4:BULK M7:DRN 0.001
R27 M4:BULK M7:BULK 0.001
R28 M4:BULK M5:BULK 0.001
R29 M4:BULK M10:BULK 0.001
R30 M4:BULK M11:BULK 0.001
R31 M4:BULK M8:BULK 0.001
R32 M4:BULK M9:BULK 0.001
R33 M4:BULK M6:BULK 0.001
R34 M4:BULK M12:BULK 0.001
R35 M4:BULK M13:BULK 0.001
R36 M4:BULK M2:BULK 0.001
R37 M4:BULK M1:BULK 0.001
R38 M4:BULK M3:BULK 0.001
R39 M12:SRC M7:DRN 8e-10
R40 M12:SRC GND 31.0176
R41 M12:SRC M13:DRN 0.001
R42 M3:DRN M7:DRN 1.875e-09
R43 M11:DRN M7:DRN 47.1809
R44 M11:DRN GND 32.2043
R45 M11:DRN M10:SRC 0.001
R46 GND M7:DRN 1.06519
R47 M7:DRN M6:DRN 0.001
R48 M15:DRN M14:SRC 81.9545
R49 M15:DRN M5:DRN 78.9176
R50 M15:DRN M2:DRN 68.8702
R51 M14:SRC M17:DRN 0.001
R52 M14:SRC M5:DRN 68.6718
R53 M14:SRC M2:DRN 78.6751
R54 M5:DRN M2:DRN 75.7597
R55 M5:DRN M4:DRN 0.001
R56 M15:GATE M16:DRN 264.942
R57 M15:GATE M13:SRC 264.526
R58 M15:GATE M1:GATE 276.219
R59 M16:DRN M13:SRC 41.0216
R60 M16:DRN M1:GATE 447.432
R61 M1:GATE M13:SRC 446.731
R62 M23:SRC Z 9.33144
R63 Z M3:SRC 9.20759
R64 N_4:1 M9:SRC 26.0503
R65 N_4:1 M19:DRN 25.3883
R66 N_4:1 M20:SRC 18.25
R67 N_4:1 M1:DRN 19.0227
R68 M19:DRN M9:SRC 125.319
R69 M19:DRN M18:DRN 0.001
R70 M9:SRC M8:DRN 0.001
R71 M26:DRN M14:DRN 53.8838
R72 M26:DRN M12:DRN 54.9942
R73 M14:DRN M12:DRN 55.7495
R74 M12:DRN M5:SRC 0.001
R75 M23:GATE M20:DRN 224.825
R76 M23:GATE M1:SRC 216.057
R77 M23:GATE M3:GATE 231.323
R78 M20:DRN M1:SRC 44.4352
R79 M20:DRN M3:GATE 207.928
R80 M20:DRN M15:SRC 0.001
R81 M3:GATE M1:SRC 199.819
R82 M1:SRC M2:SRC 0.001
R83 M26:GATE M12:GATE 305.443
R84 M26:GATE I3 93.2367
R85 I3 M12:GATE 76.4373
R86 M20:GATE M16:GATE 236.52
R87 M20:GATE S1 106.089
R88 M16:GATE M13:GATE 80.46
R89 M13:GATE M2:GATE 177.12
R90 M22:SRC M7:SRC 36.5689
R91 M22:SRC M17:SRC 0.001
R92 M7:SRC M4:SRC 0.001
R93 VDD:1 M24:SRC 2.7759
R94 VDD:1 M21:SRC 20.1294
R95 VDD:1 M26:SRC 1.89258
R96 VDD:1 M23:DRN 10.0663
R97 VDD:1 VDD 0.741753
R98 M20:BULK M24:SRC 0.001
R99 M20:BULK M21:SRC 0.00257202
R100 M20:BULK M26:SRC 0.00237417
R101 M20:BULK M26:BULK 0.001
R102 M20:BULK M15:BULK 0.001
R103 M20:BULK M25:BULK 0.001
R104 M20:BULK M22:BULK 0.001
R105 M20:BULK M16:BULK 0.001
R106 M20:BULK M24:BULK 0.001
R107 M20:BULK M21:BULK 0.001
R108 M20:BULK M19:BULK 0.001
R109 M20:BULK M23:DRN 0.00411523
R110 M20:BULK M18:BULK 0.001
R111 M20:BULK M23:BULK 0.001
R112 M20:BULK M14:BULK 0.001
R113 M20:BULK M17:BULK 0.001
R114 VDD M24:SRC 2.07113
R115 M23:DRN M26:SRC 5.03704e-10
R116 M26:SRC M16:SRC 0.001
R117 M26:SRC M24:SRC 2.1e-09
R118 M24:SRC M21:SRC 5e-10
R119 M24:SRC M25:DRN 0.001
R120 M21:SRC M22:DRN 0.001
R121 N_11:1 M9:GATE 41.1692
R122 N_11:1 M10:DRN 21.435
R123 N_11:1 M24:DRN 22.3505
R124 N_11:1 M18:GATE 66.5728
R125 N_11:1 M4:GATE 49.7667
R126 M14:GATE M4:GATE 90.72
R127 M24:DRN M10:DRN 279.849
R128 M24:DRN M18:GATE 549.502
R129 M18:GATE M10:DRN 833.554
c_1 M25:SRC 0 1.27398e-17 
c_2 M11:SRC 0 9.88483e-18 
c_3 M22:GATE 0 1.02871e-17 
c_4 I2 0 1.19998e-17 
c_5 M7:GATE 0 3.5337e-18 
c_6 M21:GATE I2 2.20098e-18 
c_7 M21:GATE M22:GATE 6.11373e-18 
c_8 M21:GATE 0 8.17751e-18 
c_9 I0 I2 5.16613e-17 
c_10 I0 M22:GATE 1.91559e-18 
c_11 I0 0 1.28505e-17 
c_12 M6:GATE I2 2.08444e-17 
c_13 M6:GATE M7:GATE 5.49641e-19 
c_14 M6:GATE 0 1.52333e-18 
c_15 M25:GATE M25:SRC 7.9422e-18 
c_16 M25:GATE 0 2.007e-18 
c_17 I1 M11:SRC 5.41947e-17 
c_18 I1 M25:SRC 1.34497e-17 
c_19 I1 0 1.22089e-18 
c_20 M11:GATE M11:SRC 1.02652e-17 
c_21 M11:GATE M25:SRC 2.71513e-18 
c_22 M11:GATE 0 3.31731e-18 
c_23 M5:GATE I2 1.00593e-19 
c_24 M5:GATE M7:GATE 4.15784e-19 
c_25 M5:GATE 0 2.38039e-19 
c_26 M24:GATE I1 2.25062e-18 
c_27 M24:GATE M25:SRC 2.93426e-20 
c_28 M24:GATE M25:GATE 7.12385e-18 
c_29 M24:GATE 0 1.49323e-18 
c_30 M17:GATE I0 1.88636e-19 
c_31 M17:GATE I2 6.12449e-19 
c_32 M17:GATE M22:GATE 6.50977e-18 
c_33 M19:GATE M11:SRC 2.19341e-17 
c_34 M19:GATE I0 1.16637e-19 
c_35 M19:GATE I2 1.08749e-19 
c_36 M19:GATE M22:GATE 1.76146e-20 
c_37 M19:GATE I1 2.4809e-18 
c_38 M19:GATE M25:SRC 2.00516e-20 
c_39 M19:GATE M11:GATE 3.35471e-18 
c_40 M19:GATE M25:GATE 1.67603e-18 
c_41 M19:GATE 0 2.37047e-17 
c_42 S0 M11:SRC 3.19868e-19 
c_43 S0 I0 1.44673e-17 
c_44 S0 I2 9.98458e-20 
c_45 S0 M22:GATE 1.8593e-17 
c_46 S0 I1 8.71505e-17 
c_47 S0 M25:SRC 6.04846e-17 
c_48 S0 M11:GATE 8.14758e-19 
c_49 S0 M25:GATE 8.75194e-18 
c_50 S0 M21:GATE 6.62045e-19 
c_51 S0 0 1.36525e-18 
c_52 M10:GATE M11:SRC 4.10128e-20 
c_53 M10:GATE M6:GATE 9.8066e-20 
c_54 M10:GATE I1 1.12967e-17 
c_55 M10:GATE M25:SRC 8.81244e-20 
c_56 M10:GATE M11:GATE 2.69703e-18 
c_57 M10:GATE 0 1.88791e-18 
c_58 M8:GATE M11:SRC 1.42565e-17 
c_59 M8:GATE M6:GATE 1.26042e-19 
c_60 M8:GATE I0 6.87262e-18 
c_61 M8:GATE I2 3.08289e-20 
c_62 M8:GATE M11:GATE 2.06237e-18 
c_63 M8:GATE 0 7.91895e-18 
c_64 M21:DRN S0 1.74223e-17 
c_65 M21:DRN M8:GATE 2.16637e-17 
c_66 M21:DRN M19:GATE 1.5929e-17 
c_67 M21:DRN M6:GATE 8.29823e-20 
c_68 M21:DRN I0 1.39068e-17 
c_69 M21:DRN 0 1.30307e-17 
c_70 M6:SRC S0 8.52115e-19 
c_71 M6:SRC M8:GATE 2.86456e-18 
c_72 M6:SRC M19:GATE 1.71576e-18 
c_73 M6:SRC M6:GATE 2.79793e-18 
c_74 M6:SRC I0 7.35644e-17 
c_75 M6:SRC 0 2.464e-17 
c_76 M4:BULK M8:GATE 2.96062e-18 
c_77 M4:BULK M19:GATE 3.02276e-19 
c_78 M4:BULK M6:GATE 8.20776e-18 
c_79 M4:BULK I0 1.96623e-19 
c_80 M4:BULK I2 2.49893e-18 
c_81 M4:BULK M10:GATE 9.24483e-18 
c_82 M4:BULK I1 2.50815e-18 
c_83 M4:BULK M25:SRC 2.53916e-18 
c_84 M4:BULK M11:GATE 1.411e-17 
c_85 M4:BULK M7:GATE 1.102e-17 
c_86 M4:BULK M5:GATE 9.50405e-18 
c_87 M4:BULK M24:GATE 5.65667e-18 
c_88 M4:BULK 0 2.60864e-18 
c_89 M12:SRC M7:GATE 8.32982e-20 
c_90 M12:SRC M5:GATE 2.65876e-19 
c_91 M12:SRC 0 9.38496e-18 
c_92 M3:DRN 0 3.02698e-17 
c_93 M11:DRN S0 1.34734e-18 
c_94 M11:DRN M8:GATE 4.77862e-20 
c_95 M11:DRN M19:GATE 1.31301e-20 
c_96 M11:DRN M10:GATE 1.46261e-17 
c_97 M11:DRN I1 1.27393e-17 
c_98 M11:DRN M25:SRC 3.59254e-19 
c_99 M11:DRN M24:GATE 7.70965e-18 
c_100 M11:DRN 0 9.01209e-18 
c_101 GND S0 4.15435e-18 
c_102 GND M11:SRC 1.2056e-18 
c_103 GND M8:GATE 2.0784e-18 
c_104 GND M19:GATE 2.31283e-20 
c_105 GND M6:GATE 4.07697e-18 
c_106 GND I0 2.37243e-18 
c_107 GND I2 2.53022e-18 
c_108 GND M10:GATE 9.19294e-18 
c_109 GND I1 2.51489e-18 
c_110 GND M25:SRC 1.1025e-18 
c_111 GND M11:GATE 5.79589e-18 
c_112 GND M7:GATE 3.78117e-18 
c_113 GND M5:GATE 2.72641e-18 
c_114 GND 0 1.70695e-16 
c_115 M7:DRN S0 2.24758e-19 
c_116 M7:DRN M11:SRC 1.24922e-17 
c_117 M7:DRN M8:GATE 4.78221e-18 
c_118 M7:DRN M19:GATE 6.01386e-20 
c_119 M7:DRN M6:GATE 2.42301e-17 
c_120 M7:DRN I0 1.54203e-17 
c_121 M7:DRN I2 2.20994e-18 
c_122 M7:DRN M10:GATE 9.18621e-18 
c_123 M7:DRN I1 3.09409e-19 
c_124 M7:DRN M11:GATE 9.42673e-18 
c_125 M7:DRN M7:GATE 2.49146e-17 
c_126 M7:DRN M17:GATE 1.52986e-20 
c_127 M7:DRN M5:GATE 5.6819e-18 
c_128 M7:DRN 0 2.54025e-16 
c_129 M15:DRN M7:DRN 1.06835e-19 
c_130 M15:DRN M5:GATE 1.06348e-17 
c_131 M15:DRN 0 7.38188e-18 
c_132 M14:SRC M7:DRN 4.13407e-20 
c_133 M14:SRC S0 2.69492e-17 
c_134 M14:SRC M17:GATE 2.7931e-18 
c_135 M14:SRC 0 7.81859e-18 
c_136 M5:DRN M7:DRN 1.66877e-17 
c_137 M5:DRN GND 1.10939e-18 
c_138 M5:DRN M17:GATE 1.20374e-17 
c_139 M5:DRN M12:SRC 5.81592e-18 
c_140 M2:DRN M7:DRN 1.05199e-17 
c_141 M2:DRN GND 1.62944e-16 
c_142 M2:DRN S0 1.39207e-18 
c_143 M2:DRN M4:BULK 7.30898e-18 
c_144 M2:DRN M17:GATE 6.4209e-18 
c_145 M2:DRN M12:SRC 1.73281e-18 
c_146 M2:DRN 0 3.16117e-18 
c_147 M15:GATE M14:SRC 7.10862e-17 
c_148 M15:GATE M4:BULK 6.48403e-18 
c_149 M15:GATE M2:DRN 2.14958e-19 
c_150 M15:GATE M3:DRN 7.59776e-19 
c_151 M15:GATE 0 8.41721e-18 
c_152 M16:DRN M7:DRN 7.93312e-20 
c_153 M16:DRN M5:DRN 1.05983e-16 
c_154 M16:DRN M15:DRN 3.50543e-17 
c_155 M16:DRN 0 1.56403e-17 
c_156 M1:GATE M7:DRN 1.35089e-17 
c_157 M1:GATE GND 6.1046e-18 
c_158 M1:GATE M4:BULK 4.27183e-18 
c_159 M1:GATE M12:SRC 8.37309e-20 
c_160 M1:GATE M2:DRN 5.76697e-20 
c_161 M1:GATE 0 2.15433e-17 
c_162 M13:SRC M7:DRN 2.17059e-18 
c_163 M13:SRC GND 3.40911e-18 
c_164 M13:SRC M4:BULK 1.07897e-17 
c_165 M13:SRC M5:DRN 5.01119e-18 
c_166 M13:SRC M15:DRN 1.83155e-17 
c_167 M13:SRC M2:DRN 1.62676e-17 
c_168 M13:SRC M3:DRN 1.51336e-20 
c_169 M13:SRC 0 1.53546e-17 
c_170 M23:SRC M7:DRN 3.34231e-20 
c_171 M23:SRC 0 6.22038e-18 
c_172 Z M7:DRN 8.58431e-19 
c_173 Z GND 4.34679e-17 
c_174 Z M4:BULK 4.78041e-19 
c_175 Z 0 5.84556e-17 
c_176 M3:SRC GND 2.11756e-18 
c_177 M3:SRC M7:DRN 1.06416e-17 
c_178 M3:SRC 0 1.99307e-18 
c_179 N_4:1 M6:SRC 3.81528e-17 
c_180 N_4:1 S0 2.06423e-16 
c_181 N_4:1 M11:SRC 4.55888e-17 
c_182 N_4:1 M8:GATE 1.83061e-17 
c_183 N_4:1 M19:GATE 2.64118e-18 
c_184 N_4:1 M21:DRN 9.23089e-17 
c_185 N_4:1 I0 3.88333e-17 
c_186 N_4:1 M14:SRC 4.30676e-17 
c_187 N_4:1 M25:SRC 1.2432e-19 
c_188 N_4:1 M17:GATE 1.35047e-17 
c_189 N_4:1 M5:GATE 3.57633e-19 
c_190 N_4:1 M16:DRN 1.43224e-18 
c_191 N_4:1 M13:SRC 2.86731e-17 
c_192 N_4:1 M15:DRN 5.09241e-17 
c_193 N_4:1 M2:DRN 3.64554e-18 
c_194 N_4:1 M1:GATE 8.29823e-20 
c_195 N_4:1 M21:GATE 7.383e-18 
c_196 N_4:1 M15:GATE 5.44772e-18 
c_197 N_4:1 0 1.66423e-17 
c_198 M20:SRC M13:SRC 8.02093e-19 
c_199 M20:SRC M15:DRN 4.27557e-19 
c_200 M20:SRC M2:DRN 1.3624e-19 
c_201 M20:SRC M15:GATE 3.48772e-20 
c_202 M20:SRC 0 1.64673e-18 
c_203 M1:DRN M13:SRC 1.03478e-17 
c_204 M1:DRN M2:DRN 1.00644e-18 
c_205 M1:DRN M1:GATE 1.91763e-17 
c_206 M1:DRN 0 4.17337e-17 
c_207 M19:DRN S0 4.03729e-18 
c_208 M19:DRN M11:SRC 7.34754e-19 
c_209 M19:DRN M8:GATE 1.26336e-17 
c_210 M19:DRN M19:GATE 2.81352e-17 
c_211 M19:DRN M21:DRN 1.34989e-18 
c_212 M19:DRN M25:SRC 6.99627e-19 
c_213 M19:DRN M5:GATE 1.02699e-17 
c_214 M9:SRC M6:SRC 7.25634e-18 
c_215 M9:SRC M11:SRC 1.01324e-18 
c_216 M9:SRC M8:GATE 2.03494e-17 
c_217 M9:SRC M19:GATE 3.80434e-18 
c_218 M9:SRC M21:DRN 2.5434e-19 
c_219 M9:SRC 0 8.11015e-18 
c_220 M26:DRN M14:SRC 3.61713e-20 
c_221 M26:DRN N_4:1 1.60907e-17 
c_222 M26:DRN M17:GATE 7.5733e-18 
c_223 M26:DRN M5:DRN 2.37888e-18 
c_224 M26:DRN M5:GATE 7.30634e-17 
c_225 M26:DRN M15:DRN 6.36904e-17 
c_226 M26:DRN 0 3.3583e-17 
c_227 M14:DRN M15:DRN 3.74185e-17 
c_228 M14:DRN M14:SRC 9.8378e-19 
c_229 M14:DRN M5:DRN 5.71257e-18 
c_230 M14:DRN M19:DRN 6.56973e-18 
c_231 M14:DRN S0 4.27595e-17 
c_232 M12:DRN M9:SRC 6.33485e-17 
c_233 M12:DRN M5:DRN 5.50506e-17 
c_234 M12:DRN M5:GATE 2.64388e-17 
c_235 M12:DRN M2:DRN 5.86552e-21 
c_236 M12:DRN 0 2.57406e-17 
c_237 M23:GATE M14:SRC 3.47234e-17 
c_238 M23:GATE M20:SRC 9.86064e-19 
c_239 M23:GATE M1:GATE 2.29925e-17 
c_240 M23:GATE M23:SRC 3.51787e-17 
c_241 M23:GATE Z 1.58829e-17 
c_242 M23:GATE 0 1.40096e-17 
c_243 M20:DRN M7:DRN 4.7354e-20 
c_244 M20:DRN M14:SRC 2.43127e-17 
c_245 M20:DRN N_4:1 1.66436e-16 
c_246 M20:DRN M16:DRN 8.17898e-18 
c_247 M20:DRN M15:DRN 8.63487e-19 
c_248 M20:DRN M20:SRC 1.30343e-18 
c_249 M20:DRN M3:SRC 9.20699e-18 
c_250 M20:DRN M23:SRC 1.74297e-19 
c_251 M20:DRN Z 8.01807e-17 
c_252 M20:DRN M15:GATE 2.41983e-17 
c_253 M20:DRN 0 4.70688e-22 
c_254 M3:GATE M7:DRN 2.40823e-17 
c_255 M3:GATE GND 5.58804e-18 
c_256 M3:GATE M14:SRC 4.07304e-17 
c_257 M3:GATE M4:BULK 2.93618e-18 
c_258 M3:GATE M1:GATE 7.96635e-19 
c_259 M3:GATE M3:SRC 2.85275e-17 
c_260 M3:GATE Z 2.76538e-17 
c_261 M1:SRC M7:DRN 1.34528e-17 
c_262 M1:SRC GND 8.62885e-17 
c_263 M1:SRC M4:BULK 1.04949e-17 
c_264 M1:SRC N_4:1 2.17697e-17 
c_265 M1:SRC M5:DRN 1.80851e-17 
c_266 M1:SRC M12:SRC 6.35719e-21 
c_267 M1:SRC M16:DRN 1.61979e-17 
c_268 M1:SRC M13:SRC 1.08514e-20 
c_269 M1:SRC M15:DRN 3.94898e-19 
c_270 M1:SRC M2:DRN 7.98099e-19 
c_271 M1:SRC M20:SRC 2.43462e-19 
c_272 M1:SRC M1:GATE 1.9683e-17 
c_273 M1:SRC M1:DRN 9.15654e-18 
c_274 M1:SRC M3:DRN 8.20305e-18 
c_275 M1:SRC M23:SRC 7.99026e-20 
c_276 M1:SRC 0 5.46672e-19 
c_277 M26:GATE S0 2.75011e-20 
c_278 M26:GATE N_4:1 9.41714e-18 
c_279 M26:GATE M17:GATE 8.18942e-18 
c_280 M26:GATE M26:DRN 1.96088e-17 
c_281 M26:GATE M16:DRN 1.19401e-19 
c_282 M26:GATE M13:SRC 1.11638e-18 
c_283 M26:GATE M15:DRN 5.20093e-18 
c_284 M26:GATE M15:GATE 5.97831e-20 
c_285 M26:GATE 0 4.34706e-18 
c_286 I3 M7:DRN 5.29574e-20 
c_287 I3 GND 9.01415e-19 
c_288 I3 M4:BULK 6.0184e-18 
c_289 I3 M14:DRN 9.1128e-17 
c_290 I3 N_4:1 1.0263e-17 
c_291 I3 M17:GATE 7.28917e-18 
c_292 I3 M5:DRN 1.26402e-17 
c_293 I3 M5:GATE 1.65446e-17 
c_294 I3 M26:DRN 4.43259e-18 
c_295 I3 M12:DRN 1.64869e-17 
c_296 I3 M12:SRC 2.74958e-18 
c_297 I3 M13:SRC 4.38998e-17 
c_298 I3 0 3.26506e-19 
c_299 M12:GATE M7:DRN 1.70977e-17 
c_300 M12:GATE GND 4.41326e-18 
c_301 M12:GATE M4:BULK 4.45422e-18 
c_302 M12:GATE M5:GATE 1.32608e-18 
c_303 M12:GATE M26:DRN 1.65965e-19 
c_304 M12:GATE M12:DRN 9.95218e-18 
c_305 M12:GATE M12:SRC 1.34609e-17 
c_306 M12:GATE M13:SRC 1.06706e-18 
c_307 M12:GATE M2:DRN 7.90801e-19 
c_308 M12:GATE M15:GATE 8.64007e-21 
c_309 M12:GATE 0 1.58005e-18 
c_310 M20:GATE M7:DRN 4.80084e-19 
c_311 M20:GATE M4:BULK 2.31441e-18 
c_312 M20:GATE N_4:1 3.97073e-17 
c_313 M20:GATE M16:DRN 4.15234e-19 
c_314 M20:GATE M13:SRC 6.80229e-19 
c_315 M20:GATE M15:DRN 7.80712e-18 
c_316 M20:GATE M2:DRN 3.33479e-19 
c_317 M20:GATE M20:DRN 2.28102e-17 
c_318 M20:GATE M1:SRC 1.3016e-17 
c_319 M20:GATE M1:DRN 2.25323e-18 
c_320 M20:GATE M26:GATE 1.9143e-19 
c_321 M20:GATE M15:GATE 7.15598e-18 
c_322 M20:GATE M23:GATE 7.15105e-19 
c_323 M20:GATE 0 4.7735e-19 
c_324 M16:GATE M7:DRN 9.72775e-20 
c_325 M16:GATE GND 2.05843e-19 
c_326 M16:GATE N_4:1 1.27904e-19 
c_327 M16:GATE M12:GATE 5.28988e-18 
c_328 M16:GATE M12:SRC 4.01727e-18 
c_329 M16:GATE I3 6.92146e-18 
c_330 M16:GATE M16:DRN 3.40362e-17 
c_331 M16:GATE M13:SRC 1.74763e-18 
c_332 M16:GATE M15:DRN 7.04604e-18 
c_333 M16:GATE M20:DRN 1.21487e-17 
c_334 M16:GATE M1:SRC 5.21273e-19 
c_335 M16:GATE M26:GATE 1.38081e-17 
c_336 M16:GATE M15:GATE 2.41205e-18 
c_337 M16:GATE M23:GATE 1.88426e-20 
c_338 M16:GATE 0 8.35825e-18 
c_339 S1 N_4:1 8.50068e-17 
c_340 S1 M16:DRN 2.42083e-17 
c_341 S1 M13:SRC 2.72629e-19 
c_342 S1 M1:SRC 8.16843e-17 
c_343 S1 M20:SRC 3.57383e-17 
c_344 S1 M1:DRN 7.80112e-18 
c_345 S1 M23:GATE 2.24649e-18 
c_346 S1 0 1.62918e-17 
c_347 M13:GATE M7:DRN 8.07954e-17 
c_348 M13:GATE GND 2.53919e-17 
c_349 M13:GATE M4:BULK 1.27491e-17 
c_350 M13:GATE M5:DRN 2.44755e-18 
c_351 M13:GATE M12:GATE 9.11205e-18 
c_352 M13:GATE I3 2.76061e-18 
c_353 M13:GATE M16:DRN 3.22512e-18 
c_354 M13:GATE M13:SRC 5.77748e-17 
c_355 M13:GATE M15:DRN 3.80457e-19 
c_356 M13:GATE M2:DRN 2.68606e-19 
c_357 M13:GATE M1:SRC 4.41203e-20 
c_358 M13:GATE M26:GATE 3.2025e-18 
c_359 M13:GATE 0 4.15744e-18 
c_360 M2:GATE M7:DRN 5.26184e-20 
c_361 M2:GATE GND 2.36731e-18 
c_362 M2:GATE M4:BULK 5.7426e-18 
c_363 M2:GATE N_4:1 6.62084e-19 
c_364 M2:GATE M5:DRN 1.71485e-17 
c_365 M2:GATE M12:GATE 4.79236e-20 
c_366 M2:GATE M12:SRC 2.67306e-17 
c_367 M2:GATE M16:DRN 7.93339e-18 
c_368 M2:GATE M13:SRC 8.96355e-18 
c_369 M2:GATE M2:DRN 3.86942e-17 
c_370 M2:GATE M20:DRN 5.134e-19 
c_371 M2:GATE M1:SRC 2.35768e-17 
c_372 M2:GATE M1:GATE 8.69165e-18 
c_373 M2:GATE M1:DRN 5.62285e-19 
c_374 M2:GATE M3:DRN 1.00529e-19 
c_375 M2:GATE M3:GATE 1.87572e-19 
c_376 M2:GATE 0 1.16712e-19 
c_377 M22:SRC M7:DRN 3.06777e-19 
c_378 M22:SRC S0 4.21602e-17 
c_379 M22:SRC I2 7.71211e-17 
c_380 M22:SRC M22:GATE 1.90548e-17 
c_381 M22:SRC M14:SRC 1.04894e-18 
c_382 M22:SRC N_4:1 5.34968e-18 
c_383 M22:SRC M5:DRN 2.61796e-19 
c_384 M22:SRC M5:GATE 4.21714e-20 
c_385 M22:SRC M15:DRN 5.6725e-17 
c_386 M22:SRC 0 1.86642e-17 
c_387 M7:SRC M7:DRN 1.54136e-17 
c_388 M7:SRC GND 3.13149e-19 
c_389 M7:SRC S0 5.54443e-18 
c_390 M7:SRC I2 1.27235e-17 
c_391 M7:SRC M22:GATE 3.1149e-18 
c_392 M7:SRC M14:SRC 6.19636e-18 
c_393 M7:SRC N_4:1 4.36418e-17 
c_394 M7:SRC M7:GATE 3.03626e-18 
c_395 M7:SRC M17:GATE 8.02113e-18 
c_396 M7:SRC M5:DRN 1.45583e-18 
c_397 M7:SRC M5:GATE 7.68668e-19 
c_398 M7:SRC M12:SRC 4.70688e-22 
c_399 M7:SRC M2:DRN 2.8576e-17 
c_400 M7:SRC 0 1.25212e-17 
c_401 VDD:1 S0 2.57647e-19 
c_402 VDD:1 M19:GATE 1.85325e-19 
c_403 VDD:1 I0 2.60215e-19 
c_404 VDD:1 M22:GATE 1.56286e-19 
c_405 VDD:1 N_4:1 8.4714e-17 
c_406 VDD:1 M17:GATE 1.65695e-18 
c_407 VDD:1 M12:GATE 7.95819e-20 
c_408 VDD:1 I3 9.15919e-19 
c_409 VDD:1 M16:GATE 3.24339e-18 
c_410 VDD:1 M20:GATE 2.81436e-18 
c_411 VDD:1 M1:SRC 7.30774e-18 
c_412 VDD:1 M20:SRC 1.26134e-18 
c_413 VDD:1 M23:SRC 1.35935e-18 
c_414 VDD:1 Z 3.70869e-17 
c_415 VDD:1 M24:GATE 1.54452e-18 
c_416 VDD:1 M25:GATE 1.33608e-18 
c_417 VDD:1 M21:GATE 8.62778e-19 
c_418 VDD:1 M26:GATE 1.43276e-18 
c_419 VDD:1 M23:GATE 8.22942e-18 
c_420 VDD:1 S1 2.53629e-17 
c_421 VDD:1 0 4.84691e-17 
c_422 M20:BULK S0 1.39263e-17 
c_423 M20:BULK M19:GATE 2.64904e-18 
c_424 M20:BULK M6:GATE 3.41136e-18 
c_425 M20:BULK I0 1.6607e-18 
c_426 M20:BULK I2 8.61797e-19 
c_427 M20:BULK M22:GATE 3.717e-18 
c_428 M20:BULK N_4:1 2.28664e-17 
c_429 M20:BULK M10:GATE 3.25647e-18 
c_430 M20:BULK M19:DRN 1.91308e-18 
c_431 M20:BULK M7:GATE 3.49608e-18 
c_432 M20:BULK M17:GATE 2.59716e-17 
c_433 M20:BULK M5:GATE 1.96462e-18 
c_434 M20:BULK I3 1.67883e-18 
c_435 M20:BULK M16:GATE 9.39165e-18 
c_436 M20:BULK M20:DRN 2.35042e-18 
c_437 M20:BULK M20:GATE 1.9386e-17 
c_438 M20:BULK M1:SRC 5.47869e-18 
c_439 M20:BULK M23:SRC 6.22358e-18 
c_440 M20:BULK Z 6.36266e-18 
c_441 M20:BULK M24:GATE 6.27495e-18 
c_442 M20:BULK M25:GATE 1.0794e-17 
c_443 M20:BULK M21:GATE 4.07389e-18 
c_444 M20:BULK M26:GATE 7.87782e-18 
c_445 M20:BULK M23:GATE 3.67247e-18 
c_446 M20:BULK S1 1.33277e-18 
c_447 M20:BULK 0 6.00262e-18 
c_448 VDD S0 2.33004e-16 
c_449 VDD I0 2.37673e-19 
c_450 VDD M22:GATE 4.20088e-18 
c_451 VDD N_4:1 1.67183e-16 
c_452 VDD M16:GATE 3.56501e-18 
c_453 VDD M20:DRN 9.76574e-19 
c_454 VDD M20:GATE 3.10995e-17 
c_455 VDD M1:SRC 1.29129e-18 
c_456 VDD M20:SRC 5.36693e-20 
c_457 VDD M23:SRC 2.10925e-18 
c_458 VDD Z 2.96914e-17 
c_459 VDD M24:GATE 5.45046e-18 
c_460 VDD M25:GATE 4.19228e-18 
c_461 VDD M21:GATE 3.36912e-18 
c_462 VDD M26:GATE 4.79389e-18 
c_463 VDD M23:GATE 5.91801e-18 
c_464 VDD S1 4.49526e-19 
c_465 VDD 0 1.77159e-16 
c_466 M23:DRN N_4:1 2.33404e-18 
c_467 M23:DRN M16:GATE 3.72075e-18 
c_468 M23:DRN M20:DRN 6.09841e-18 
c_469 M23:DRN M20:GATE 1.03168e-17 
c_470 M23:DRN M20:SRC 3.2925e-17 
c_471 M23:DRN M23:SRC 9.859e-19 
c_472 M23:DRN Z 4.47704e-19 
c_473 M23:DRN M23:GATE 4.54853e-17 
c_474 M23:DRN S1 1.01173e-18 
c_475 M23:DRN 0 7.44553e-18 
c_476 M26:SRC S0 8.84037e-19 
c_477 M26:SRC M22:GATE 5.20109e-22 
c_478 M26:SRC N_4:1 7.73144e-18 
c_479 M26:SRC M12:GATE 2.82854e-18 
c_480 M26:SRC I3 3.14194e-18 
c_481 M26:SRC M16:GATE 4.19837e-17 
c_482 M26:SRC M20:DRN 8.2633e-20 
c_483 M26:SRC M20:GATE 4.21266e-17 
c_484 M26:SRC M1:SRC 9.61521e-21 
c_485 M26:SRC M20:SRC 4.10883e-20 
c_486 M26:SRC M1:DRN 1.06049e-22 
c_487 M26:SRC M23:SRC 7.58727e-19 
c_488 M26:SRC Z 8.5269e-19 
c_489 M26:SRC M26:GATE 2.0186e-17 
c_490 M26:SRC M23:GATE 5.15617e-18 
c_491 M26:SRC S1 9.1308e-20 
c_492 M26:SRC 0 2.81499e-17 
c_493 M24:SRC M9:SRC 8.7017e-20 
c_494 M24:SRC S0 8.33996e-17 
c_495 M24:SRC M19:GATE 5.58971e-19 
c_496 M24:SRC I0 3.1418e-19 
c_497 M24:SRC I2 1.19314e-19 
c_498 M24:SRC M22:GATE 9.49751e-18 
c_499 M24:SRC N_4:1 1.60505e-18 
c_500 M24:SRC I1 1.5917e-18 
c_501 M24:SRC M19:DRN 3.15155e-18 
c_502 M24:SRC M5:GATE 2.53229e-19 
c_503 M24:SRC I3 6.80906e-20 
c_504 M24:SRC M16:GATE 1.59493e-18 
c_505 M24:SRC M20:DRN 5.23863e-18 
c_506 M24:SRC M20:GATE 3.34653e-17 
c_507 M24:SRC M1:SRC 6.15775e-20 
c_508 M24:SRC M20:SRC 7.79917e-18 
c_509 M24:SRC M1:DRN 8.33668e-20 
c_510 M24:SRC M3:SRC 2.8543e-20 
c_511 M24:SRC M23:SRC 6.40372e-18 
c_512 M24:SRC Z 1.37762e-19 
c_513 M24:SRC M24:GATE 3.10783e-17 
c_514 M24:SRC M25:GATE 3.05385e-17 
c_515 M24:SRC M21:GATE 9.3648e-18 
c_516 M24:SRC M26:GATE 7.17582e-18 
c_517 M24:SRC M23:GATE 4.35799e-18 
c_518 M24:SRC 0 2.12308e-16 
c_519 M21:SRC S0 7.59441e-18 
c_520 M21:SRC I0 9.39719e-18 
c_521 M21:SRC I2 3.33006e-18 
c_522 M21:SRC M22:GATE 1.86708e-17 
c_523 M21:SRC N_4:1 6.58473e-18 
c_524 M21:SRC M19:DRN 3.47244e-20 
c_525 M21:SRC M20:GATE 1.06049e-22 
c_526 M21:SRC Z 5.11622e-20 
c_527 M21:SRC M25:GATE 2.96445e-19 
c_528 M21:SRC M21:GATE 1.91535e-17 
c_529 M21:SRC M26:GATE 5.20109e-22 
c_530 M21:SRC 0 6.78289e-18 
c_531 N_11:1 M7:DRN 1.09072e-17 
c_532 N_11:1 M6:SRC 1.93374e-17 
c_533 N_11:1 M9:SRC 2.42332e-17 
c_534 N_11:1 GND 3.02066e-16 
c_535 N_11:1 M24:SRC 1.55644e-17 
c_536 N_11:1 S0 1.59763e-16 
c_537 N_11:1 M11:DRN 5.24248e-18 
c_538 N_11:1 M11:SRC 9.32765e-18 
c_539 N_11:1 M8:GATE 2.11989e-18 
c_540 N_11:1 M19:GATE 1.68384e-17 
c_541 N_11:1 M6:GATE 5.50904e-18 
c_542 N_11:1 M21:DRN 2.81842e-17 
c_543 N_11:1 I0 1.27356e-17 
c_544 N_11:1 M22:GATE 6.2172e-18 
c_545 N_11:1 M7:SRC 6.22403e-17 
c_546 N_11:1 M22:SRC 2.71969e-18 
c_547 N_11:1 M14:SRC 1.87686e-17 
c_548 N_11:1 M4:BULK 1.46353e-17 
c_549 N_11:1 N_4:1 1.20859e-18 
c_550 N_11:1 M10:GATE 1.76579e-19 
c_551 N_11:1 I1 3.49936e-17 
c_552 N_11:1 M25:SRC 1.0053e-16 
c_553 N_11:1 M11:GATE 4.6528e-19 
c_554 N_11:1 M19:DRN 4.39007e-17 
c_555 N_11:1 M21:SRC 1.27253e-19 
c_556 N_11:1 M7:GATE 1.31943e-18 
c_557 N_11:1 M17:GATE 4.63899e-17 
c_558 N_11:1 M5:DRN 1.73691e-17 
c_559 N_11:1 M5:GATE 1.91434e-17 
c_560 N_11:1 M12:DRN 5.82656e-19 
c_561 N_11:1 M23:DRN 2.24766e-19 
c_562 N_11:1 VDD 1.42056e-16 
c_563 N_11:1 M24:GATE 1.34141e-17 
c_564 N_11:1 M25:GATE 1.91757e-17 
c_565 N_11:1 M21:GATE 7.14478e-18 
c_566 N_11:1 VDD:1 1.6275e-20 
c_567 N_11:1 0 2.93221e-18 
c_568 M14:GATE M6:SRC 1.17373e-19 
c_569 M14:GATE M24:SRC 1.37408e-18 
c_570 M14:GATE S0 1.67237e-17 
c_571 M14:GATE M6:GATE 2.47088e-20 
c_572 M14:GATE I0 6.54328e-20 
c_573 M14:GATE I2 1.67759e-18 
c_574 M14:GATE M22:GATE 9.0657e-19 
c_575 M14:GATE M22:SRC 3.5805e-18 
c_576 M14:GATE M14:SRC 1.88794e-17 
c_577 M14:GATE M4:BULK 6.86302e-18 
c_578 M14:GATE M14:DRN 1.4774e-17 
c_579 M14:GATE N_4:1 5.06959e-20 
c_580 M14:GATE M20:BULK 9.41412e-18 
c_581 M14:GATE M19:DRN 7.20724e-18 
c_582 M14:GATE M7:GATE 5.94813e-19 
c_583 M14:GATE M17:GATE 1.08826e-17 
c_584 M14:GATE M26:DRN 5.4051e-18 
c_585 M14:GATE M12:DRN 5.99126e-21 
c_586 M14:GATE M2:DRN 1.0089e-17 
c_587 M14:GATE VDD 1.21886e-18 
c_588 M14:GATE 0 2.32286e-18 
c_589 M4:GATE M7:DRN 8.46762e-21 
c_590 M4:GATE S0 3.71453e-18 
c_591 M4:GATE M6:GATE 2.94485e-21 
c_592 M4:GATE I2 1.62656e-19 
c_593 M4:GATE M7:SRC 1.42549e-17 
c_594 M4:GATE M22:SRC 2.05745e-18 
c_595 M4:GATE M5:DRN 1.77835e-17 
c_596 M4:GATE M5:GATE 7.8432e-18 
c_597 M4:GATE M2:DRN 3.53879e-18 
c_598 M4:GATE 0 1.04518e-18 
c_599 M24:DRN M7:DRN 1.30159e-17 
c_600 M24:DRN GND 5.08436e-17 
c_601 M24:DRN M24:SRC 9.19407e-18 
c_602 M24:DRN S0 2.46208e-19 
c_603 M24:DRN M20:BULK 2.73182e-18 
c_604 M24:DRN M25:SRC 1.18748e-18 
c_605 M24:DRN VDD 1.98178e-18 
c_606 M24:DRN M24:GATE 1.68548e-17 
c_607 M24:DRN M25:GATE 7.74427e-20 
c_608 M24:DRN 0 9.42367e-18 
c_609 M18:GATE M7:DRN 1.76906e-20 
c_610 M18:GATE GND 1.23548e-20 
c_611 M18:GATE M24:SRC 2.34682e-18 
c_612 M18:GATE S0 1.23251e-17 
c_613 M18:GATE M11:SRC 4.29415e-18 
c_614 M18:GATE M19:GATE 9.45539e-18 
c_615 M18:GATE M21:DRN 5.60099e-19 
c_616 M18:GATE I0 1.09592e-19 
c_617 M18:GATE N_4:1 3.31648e-18 
c_618 M18:GATE M20:BULK 3.57471e-18 
c_619 M18:GATE I1 7.16024e-19 
c_620 M18:GATE M25:SRC 7.79138e-18 
c_621 M18:GATE M19:DRN 5.42408e-18 
c_622 M18:GATE M24:GATE 9.40432e-20 
c_623 M18:GATE M25:GATE 2.92617e-18 
c_624 M18:GATE VDD:1 3.46693e-19 
c_625 M18:GATE 0 3.87015e-17 
c_626 M9:GATE M7:DRN 7.75597e-18 
c_627 M9:GATE M6:SRC 1.87408e-17 
c_628 M9:GATE M9:SRC 1.68649e-17 
c_629 M9:GATE GND 3.7634e-18 
c_630 M9:GATE S0 4.23655e-22 
c_631 M9:GATE M11:SRC 7.13575e-19 
c_632 M9:GATE M8:GATE 1.34482e-17 
c_633 M9:GATE M19:GATE 5.07906e-18 
c_634 M9:GATE M21:DRN 4.94154e-21 
c_635 M9:GATE I0 5.84011e-18 
c_636 M9:GATE I2 2.93367e-19 
c_637 M9:GATE M4:BULK 6.01969e-18 
c_638 M9:GATE N_4:1 7.27522e-18 
c_639 M9:GATE I1 4.66901e-20 
c_640 M9:GATE M11:GATE 6.73417e-20 
c_641 M9:GATE M19:DRN 6.97313e-19 
c_642 M9:GATE 0 5.38865e-18 
c_643 M10:DRN M7:DRN 9.88443e-18 
c_644 M10:DRN GND 1.61644e-18 
c_645 M10:DRN M24:SRC 4.36823e-20 
c_646 M10:DRN S0 1.68212e-17 
c_647 M10:DRN M11:DRN 7.64805e-19 
c_648 M10:DRN M11:SRC 7.35905e-19 
c_649 M10:DRN I2 3.7555e-17 
c_650 M10:DRN M20:BULK 1.0706e-17 
c_651 M10:DRN I1 1.12778e-20 
c_652 M10:DRN 0 8.02804e-18 

.ENDS
