
.subckt INVD1  I ZN
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.15471p as=0.12636p l=0.09u nrd=0.531 nrs=0.433 pd=1.944u ps=1.548u sa=2.34e-07 sb=2.34e-07 w=0.54u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK pch ad=0.19683p as=0.16848p l=0.09u nrd=0.38 nrs=0.325 pd=2.304u ps=1.908u sa=2.34e-07 sb=2.34e-07 w=0.72u 
R1 M1:BULK M1:DRN 0.001
R2 GND M1:DRN 3.68929
R3 M2:SRC ZN 9.31289
R4 ZN M1:SRC 9.19853
R5 M2:GATE I 91.9015
R6 M2:GATE M1:GATE 289.649
R7 I M1:GATE 74.8827
R8 M2:DRN M2:BULK 0.001
R9 M2:DRN VDD 3.64463
c_1 GND 0 7.27105e-17 
c_2 M1:DRN 0 3.27954e-17 
c_3 M2:SRC M1:DRN 3.55798e-20 
c_4 M2:SRC 0 5.3518e-18 
c_5 ZN GND 7.81317e-17 
c_6 ZN M1:DRN 1.57007e-18 
c_7 ZN M1:BULK 8.13807e-18 
c_8 ZN 0 4.74243e-17 
c_9 M1:SRC M1:DRN 1.21324e-17 
c_10 M1:SRC GND 3.30943e-18 
c_11 M1:SRC 0 2.20695e-18 
c_12 M2:GATE M2:SRC 3.34781e-17 
c_13 M2:GATE ZN 9.49021e-18 
c_14 M2:GATE 0 2.06032e-17 
c_15 I M1:SRC 4.15145e-19 
c_16 I GND 2.7489e-17 
c_17 I M1:DRN 4.35576e-17 
c_18 I M1:BULK 1.34343e-17 
c_19 I ZN 7.19681e-17 
c_20 I M2:SRC 1.75822e-19 
c_21 I 0 8.93274e-18 
c_22 M1:GATE M1:BULK 3.89334e-18 
c_23 M1:GATE ZN 6.50672e-18 
c_24 M1:GATE GND 1.41074e-17 
c_25 M1:GATE M1:DRN 2.02535e-17 
c_26 M1:GATE M1:SRC 3.32033e-17 
c_27 M1:GATE 0 3.00173e-20 
c_28 M2:DRN M2:GATE 5.37986e-17 
c_29 M2:DRN M2:SRC 1.09724e-17 
c_30 M2:DRN I 1.30646e-17 
c_31 M2:DRN ZN 1.52959e-18 
c_32 M2:DRN M1:SRC 3.06117e-20 
c_33 M2:DRN 0 3.0117e-17 
c_34 M2:BULK M2:GATE 7.26033e-18 
c_35 M2:BULK M2:SRC 2.00795e-18 
c_36 M2:BULK I 1.0221e-17 
c_37 M2:BULK ZN 1.13261e-17 
c_38 VDD M2:GATE 1.30341e-17 
c_39 VDD M2:SRC 3.20151e-18 
c_40 VDD I 3.66077e-17 
c_41 VDD ZN 6.95361e-17 
c_42 VDD 0 7.61475e-17 

.ENDS
