
.subckt CKLNQD4  TE E CP Q
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.02754p as=0.0162p l=0.09u nrd=0.855 nrs=0.5 pd=0.5472u ps=0.36u sa=1.458e-06 sb=4.86e-07 w=0.18u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.0162p as=0.02916p l=0.09u nrd=0.5 nrs=0.9 pd=0.36u ps=0.4257u sa=1.188e-06 sb=7.56e-07 w=0.18u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK nch ad=0.03159p as=0.07857p l=0.09u nrd=0.433 nrs=1.078 pd=0.504u ps=1.008u sa=1.098e-06 sb=8.91e-07 w=0.27u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK nch ad=0.06642p as=0.06075p l=0.09u nrd=0.909 nrs=0.833 pd=1.062u ps=0.99u sa=4.86e-07 sb=2.25e-07 w=0.27u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.02025p as=0.05589p l=0.09u nrd=0.283 nrs=0.767 pd=0.423u ps=0.954u sa=2.07e-07 sb=1.782e-06 w=0.27u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.05589p as=0.03159p l=0.09u nrd=0.767 nrs=0.433 pd=0.954u ps=0.504u sa=1.782e-06 sb=2.07e-07 w=0.27u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.04374p as=0.04536p l=0.09u nrd=0.338 nrs=0.348 pd=0.603u ps=0.774u sa=4.86e-07 sb=7.974e-07 w=0.36u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.05589p as=0.04131p l=0.09u nrd=0.767 nrs=0.57 pd=0.954u ps=0.8208u sa=4.23e-07 sb=2.07e-07 w=0.27u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.03159p as=0.07857p l=0.09u nrd=0.433 nrs=1.078 pd=0.504u ps=1.008u sa=1.458e-06 sb=5.31e-07 w=0.27u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK nch ad=0.05589p as=0.06642p l=0.09u nrd=0.767 nrs=0.909 pd=0.954u ps=1.062u sa=2.07e-07 sb=5.04e-07 w=0.27u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.03159p as=0.02025p l=0.09u nrd=0.433 nrs=0.283 pd=0.504u ps=0.423u sa=4.5e-07 sb=1.539e-06 w=0.27u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.03159p as=0.03159p l=0.09u nrd=0.433 nrs=0.433 pd=0.504u ps=0.504u sa=7.74e-07 sb=1.215e-06 w=0.27u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.04374p as=0.05832p l=0.09u nrd=0.338 nrs=0.45 pd=0.603u ps=0.8523u sa=8.19e-07 sb=3.699e-07 w=0.36u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.04536p as=0.07452p l=0.09u nrd=0.348 nrs=0.575 pd=0.774u ps=1.134u sa=2.07e-07 sb=1.1187e-06 w=0.36u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK pch ad=0.08424p as=0.11502p l=0.09u nrd=0.162 nrs=0.222 pd=0.954u ps=1.188u sa=1.2384e-06 sb=5.31e-07 w=0.72u 
MM23 M23:DRN M23:GATE M23:SRC M23:BULK pch ad=0.08424p as=0.11016p l=0.09u nrd=0.162 nrs=0.213 pd=0.954u ps=1.3554u sa=4.329e-07 sb=1.215e-06 w=0.72u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK pch ad=0.07128p as=0.06642p l=0.09u nrd=0.549 nrs=0.51 pd=1.134u ps=0.927u sa=5.31e-07 sb=1.953e-07 w=0.36u 
MM25 M25:DRN M25:GATE M25:SRC M25:BULK pch ad=0.05913p as=0.1215p l=0.09u nrd=0.232 nrs=0.477 pd=0.738u ps=1.854u sa=1.683e-07 sb=1.863e-06 w=0.504u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK pch ad=0.07452p as=0.10125p l=0.09u nrd=0.575 nrs=0.779 pd=1.134u ps=1.4283u sa=3.384e-07 sb=2.07e-07 w=0.36u 
MM27 M27:DRN M27:GATE M27:SRC M27:BULK pch ad=0.0648p as=0.0648p l=0.09u nrd=0.125 nrs=0.125 pd=0.9u ps=0.9u sa=4.77e-07 sb=5.859e-07 w=0.72u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK pch ad=0.14904p as=0.08424p l=0.09u nrd=0.287 nrs=0.162 pd=1.854u ps=0.954u sa=1.5786e-06 sb=2.07e-07 w=0.72u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK pch ad=0.11502p as=0.08424p l=0.09u nrd=0.222 nrs=0.162 pd=1.188u ps=0.954u sa=8.415e-07 sb=8.91e-07 w=0.72u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK pch ad=0.07452p as=0.06642p l=0.09u nrd=0.575 nrs=0.51 pd=1.134u ps=0.927u sa=2.07e-07 sb=5.202e-07 w=0.36u 
MM24 M24:DRN M24:GATE M24:SRC M24:BULK pch ad=0.07695p as=0.05913p l=0.09u nrd=0.304 nrs=0.232 pd=0.9486u ps=0.738u sa=4.932e-07 sb=1.539e-06 w=0.504u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK pch ad=0.0162p as=0.0324p l=0.09u nrd=0.5 nrs=1.01 pd=0.36u ps=0.3924u sa=1.098e-06 sb=7.83e-07 w=0.18u 
MM26 M26:DRN M26:GATE M26:SRC M26:BULK pch ad=0.13122p as=0.0648p l=0.09u nrd=0.252 nrs=0.125 pd=1.5696u ps=0.9u sa=7.47e-07 sb=2.79e-07 w=0.72u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK pch ad=0.0162p as=0.05022p l=0.09u nrd=0.5 nrs=1.558 pd=0.36u ps=0.7137u sa=1.368e-06 sb=5.13e-07 w=0.18u 
MM28 M28:DRN M28:GATE M28:SRC M28:BULK pch ad=0.0648p as=0.14904p l=0.09u nrd=0.125 nrs=0.287 pd=0.9u ps=1.854u sa=2.07e-07 sb=8.793e-07 w=0.72u 
R1 M9:SRC M10:DRN 0.001
R2 M5:DRN M6:DRN 0.001
R3 M5:DRN M7:SRC 36.3527
R4 M19:DRN M17:DRN 0.001
R5 M26:DRN M8:GATE 161.053
R6 M26:DRN M5:SRC 45.6045
R7 M26:DRN M18:GATE 269.484
R8 M26:DRN M17:SRC 0.001
R9 M18:GATE M8:GATE 202.375
R10 M18:GATE M5:SRC 255.218
R11 M8:GATE M5:SRC 152.527
R12 M5:SRC M10:SRC 0.001
R13 M26:GATE M10:GATE 476.996
R14 M26:GATE M13:DRN 199.611
R15 M26:GATE M15:DRN 191.376
R16 M15:DRN M10:GATE 126.993
R17 M15:DRN M13:DRN 48.1214
R18 M13:DRN M10:GATE 132.457
R19 M27:GATE TE 98.9729
R20 M27:GATE M6:GATE 352.195
R21 TE M6:GATE 81.0215
R22 M28:GATE E 88.3007
R23 M28:GATE M7:GATE 313.066
R24 E M7:GATE 82.1343
R25 M1:SRC M2:DRN 0.001
R26 M27:SRC M28:DRN 0.001
R27 M26:SRC M27:DRN 0.001
R28 M16:DRN M15:GATE 256.23
R29 M16:DRN M13:GATE 147.228
R30 M16:DRN M14:SRC 45.72
R31 M14:SRC M15:GATE 254.588
R32 M14:SRC M13:GATE 146.284
R33 M17:GATE M15:GATE 274.32
R34 M17:GATE M5:GATE 122.04
R35 M15:GATE M13:GATE 183.485
R36 Q M12:DRN 18.2144
R37 Q M4:SRC 18.2037
R38 Q M23:DRN 9.33947
R39 Q M21:DRN 9.37491
R40 M21:DRN M23:DRN 645.353
R41 M21:DRN M20:SRC 0.001
R42 M23:DRN M22:SRC 0.001
R43 M4:SRC M11:DRN 0.001
R44 M12:DRN M3:SRC 0.001
R45 GND:1 M6:SRC 19.7416
R46 GND:1 M9:DRN 1.38021
R47 GND:1 GND 0.693802
R48 GND:1 M4:DRN 19.3179
R49 GND:1 M3:DRN 18.5572
R50 M11:SRC M12:SRC 3.96713e-10
R51 M14:BULK M6:SRC 1.05979e-05
R52 M14:BULK M9:DRN 0.00108295
R53 M14:BULK M5:BULK 0.001
R54 M14:BULK M6:BULK 0.001
R55 M14:BULK M7:BULK 0.001
R56 M14:BULK M10:BULK 0.001
R57 M14:BULK M9:BULK 0.001
R58 M14:BULK M8:BULK 0.001
R59 M14:BULK M13:BULK 0.001
R60 M14:BULK M2:BULK 0.001
R61 M14:BULK M1:BULK 0.001
R62 M14:BULK M3:BULK 0.001
R63 M14:BULK M12:BULK 0.001
R64 M14:BULK M11:BULK 0.001
R65 M14:BULK M4:BULK 0.001
R66 M14:DRN M9:DRN 2.76768e-09
R67 M14:DRN M13:SRC 0.001
R68 M3:DRN M1:DRN 0.001
R69 M12:SRC M9:DRN 1.14778e-09
R70 M4:DRN M9:DRN 491.235
R71 M6:SRC M9:DRN 1.58989e-09
R72 M6:SRC GND 3.76421
R73 M6:SRC M7:DRN 0.001
R74 GND M9:DRN 6.16102
R75 M9:DRN M8:SRC 0.001
R76 N_5:1 M8:DRN 18
R77 N_5:1 M19:GATE 52.629
R78 N_5:1 M9:GATE 128.78
R79 N_5:1 M18:DRN 18.9729
R80 N_5:1 M1:GATE 103.102
R81 N_5:1 M24:GATE 72.3034
R82 M24:GATE M1:GATE 258.9
R83 M18:DRN M19:GATE 1798.97
R84 M19:GATE M9:GATE 238.758
R85 CP:1 M16:GATE 216.306
R86 CP:1 M14:GATE 117.985
R87 CP:1 M2:GATE 38.88
R88 CP:1 CP 24.751
R89 CP:1 M25:GATE 81
R90 CP M16:GATE 440.623
R91 CP M14:GATE 240.34
R92 M14:GATE M16:GATE 216.554
R93 N_13:1 M2:SRC 51.0739
R94 N_13:1 M24:SRC 48.7388
R95 N_13:1 M3:GATE 33.6533
R96 N_13:1 M12:GATE 106.451
R97 N_13:1 N_13:2 44.2624
R98 N_13:1 M22:GATE 178.377
R99 N_13:1 M23:GATE 66.96
R100 N_13:2 M12:GATE 106.451
R101 N_13:2 M11:GATE 39.96
R102 N_13:2 M4:GATE 63.8379
R103 N_13:2 M20:GATE 106.972
R104 N_13:2 M22:GATE 178.377
R105 N_13:2 M21:GATE 66.96
R106 M22:GATE M12:GATE 428.998
R107 M20:GATE M4:GATE 285.852
R108 M24:SRC M2:SRC 58.4483
R109 M24:SRC M25:DRN 0.001
R110 VDD:1 M19:SRC 18.4139
R111 VDD:1 M16:SRC 2.99083
R112 VDD:1 M25:SRC 4.38273
R113 VDD:1 VDD:2 0.222717
R114 VDD:1 VDD 0.528228
R115 VDD:2 M25:SRC 3.09871
R116 VDD:2 M24:DRN 18.4803
R117 VDD:2 M22:DRN 18
R118 VDD:2 M20:DRN 9.54819
R119 M25:BULK M16:SRC 1.04715e-05
R120 M25:BULK M25:SRC 0.00308642
R121 M25:BULK M24:DRN 0.00385802
R122 M25:BULK M22:DRN 0.00308642
R123 M25:BULK M28:BULK 0.001
R124 M25:BULK M27:BULK 0.001
R125 M25:BULK M26:BULK 0.001
R126 M25:BULK M17:BULK 0.001
R127 M25:BULK M19:BULK 0.001
R128 M25:BULK M18:BULK 0.001
R129 M25:BULK M15:BULK 0.001
R130 M25:BULK M16:BULK 0.001
R131 M25:BULK M24:BULK 0.001
R132 M25:BULK M23:BULK 0.001
R133 M25:BULK M22:BULK 0.001
R134 M25:BULK M21:BULK 0.001
R135 M25:BULK M20:BULK 0.001
R136 VDD M16:SRC 2.75211
R137 VDD M28:SRC 9.1167
R138 M16:SRC M25:SRC 1.35e-09
R139 M16:SRC M15:SRC 0.001
R140 M22:DRN M25:SRC 5.34783e-10
R141 M22:DRN M21:SRC 0.001
R142 M25:SRC M24:DRN 5.25e-10
R143 M25:SRC M20:DRN 799.61
R144 M24:DRN M23:SRC 1.23077e-09
R145 M19:SRC M18:SRC 0.001
c_1 M9:SRC 0 2.43622e-19 
c_2 M5:DRN 0 2.68164e-19 
c_3 M7:SRC 0 1.6119e-17 
c_4 M19:DRN M9:SRC 2.24758e-19 
c_5 M26:DRN 0 1.60689e-19 
c_6 M17:SRC 0 5.78741e-20 
c_7 M18:GATE 0 1.80379e-17 
c_8 M8:GATE M9:SRC 1.82283e-18 
c_9 M8:GATE 0 1.90741e-18 
c_10 M5:SRC M5:DRN 1.6677e-18 
c_11 M5:SRC M7:SRC 3.88665e-17 
c_12 M5:SRC 0 6.07619e-18 
c_13 M26:GATE M5:SRC 3.10256e-18 
c_14 M26:GATE M18:GATE 4.80504e-21 
c_15 M26:GATE M26:DRN 1.67572e-17 
c_16 M26:GATE 0 1.14928e-17 
c_17 M15:DRN M5:DRN 4.4926e-18 
c_18 M15:DRN M19:DRN 1.47643e-18 
c_19 M15:DRN M5:SRC 1.13014e-16 
c_20 M15:DRN M18:GATE 4.0488e-18 
c_21 M15:DRN M17:SRC 3.15294e-18 
c_22 M15:DRN M7:SRC 7.03857e-18 
c_23 M15:DRN 0 9.63566e-18 
c_24 M13:DRN M9:SRC 1.81811e-19 
c_25 M13:DRN M5:DRN 2.3442e-22 
c_26 M13:DRN M8:GATE 6.9686e-18 
c_27 M13:DRN M5:SRC 4.1913e-20 
c_28 M13:DRN M26:DRN 1.70872e-16 
c_29 M13:DRN 0 5.364e-18 
c_30 M10:GATE M9:SRC 3.40288e-18 
c_31 M10:GATE M5:DRN 6.14461e-20 
c_32 M10:GATE M19:DRN 2.71339e-18 
c_33 M10:GATE M8:GATE 4.67564e-18 
c_34 M10:GATE M18:GATE 1.10287e-17 
c_35 M10:GATE M26:DRN 9.45041e-18 
c_36 M10:GATE 0 4.13208e-17 
c_37 M27:GATE M15:DRN 1.7145e-17 
c_38 M27:GATE M26:GATE 2.35588e-17 
c_39 M27:GATE 0 5.96729e-18 
c_40 TE M5:DRN 1.85772e-17 
c_41 TE M10:GATE 2.53558e-19 
c_42 TE M15:DRN 6.75644e-17 
c_43 TE M7:SRC 2.51694e-17 
c_44 TE M26:GATE 5.76512e-20 
c_45 TE 0 8.18021e-18 
c_46 M6:GATE M15:DRN 9.85604e-18 
c_47 M6:GATE M7:SRC 8.63277e-18 
c_48 M6:GATE M10:GATE 1.79779e-19 
c_49 M6:GATE 0 1.43157e-17 
c_50 M28:GATE M27:GATE 2.41678e-17 
c_51 M28:GATE TE 6.56022e-18 
c_52 M28:GATE 0 2.15306e-17 
c_53 E M5:DRN 3.14079e-17 
c_54 E M7:SRC 1.33397e-17 
c_55 E TE 1.00519e-16 
c_56 E 0 8.25164e-18 
c_57 M7:GATE M6:GATE 1.16164e-17 
c_58 M7:GATE M5:DRN 2.25786e-19 
c_59 M7:GATE M7:SRC 1.33948e-17 
c_60 M7:GATE 0 6.9948e-18 
c_61 M27:SRC TE 4.46929e-18 
c_62 M27:SRC M7:SRC 6.26307e-19 
c_63 M27:SRC 0 5.78741e-20 
c_64 M26:SRC M15:DRN 1.10376e-17 
c_65 M26:SRC M5:DRN 1.28909e-18 
c_66 M26:SRC 0 6.81677e-19 
c_67 M16:DRN M13:DRN 1.68116e-17 
c_68 M16:DRN M15:DRN 6.14631e-19 
c_69 M14:SRC M8:GATE 1.22554e-18 
c_70 M14:SRC M13:DRN 2.12394e-19 
c_71 M14:SRC M18:GATE 2.15145e-18 
c_72 M14:SRC M15:DRN 1.15829e-17 
c_73 M14:SRC M26:GATE 6.81691e-17 
c_74 M14:SRC 0 2.17028e-20 
c_75 M17:GATE M5:DRN 1.48268e-17 
c_76 M17:GATE M10:GATE 4.75623e-19 
c_77 M17:GATE M19:DRN 1.88625e-18 
c_78 M17:GATE M13:DRN 2.25163e-20 
c_79 M17:GATE M5:SRC 7.05918e-18 
c_80 M17:GATE M18:GATE 2.47526e-18 
c_81 M17:GATE M15:DRN 9.90593e-18 
c_82 M17:GATE M17:SRC 2.61726e-17 
c_83 M17:GATE M7:SRC 4.02428e-18 
c_84 M17:GATE M26:GATE 2.365e-17 
c_85 M17:GATE M26:DRN 1.42388e-17 
c_86 M17:GATE 0 1.24803e-17 
c_87 M15:GATE M10:GATE 1.39257e-17 
c_88 M15:GATE M13:DRN 1.18524e-20 
c_89 M15:GATE M18:GATE 1.0656e-18 
c_90 M15:GATE M15:DRN 2.49727e-17 
c_91 M15:GATE M26:GATE 4.01017e-20 
c_92 M15:GATE 0 1.12226e-17 
c_93 M13:GATE M8:GATE 5.52245e-20 
c_94 M13:GATE M13:DRN 6.57222e-18 
c_95 M13:GATE 0 7.76324e-18 
c_96 M5:GATE M10:GATE 1.2797e-17 
c_97 M5:GATE M5:SRC 5.0914e-17 
c_98 M5:GATE M18:GATE 3.42953e-19 
c_99 M5:GATE M15:DRN 1.90595e-17 
c_100 M5:GATE 0 1.02194e-17 
c_101 Q 0 5.44155e-18 
c_102 M21:DRN 0 3.91468e-18 
c_103 M23:DRN 0 4.27968e-18 
c_104 M4:SRC 0 1.36624e-18 
c_105 M12:DRN 0 1.38599e-18 
c_106 GND:1 M9:SRC 1.20777e-19 
c_107 GND:1 M5:DRN 6.40462e-17 
c_108 GND:1 M8:GATE 4.20133e-18 
c_109 GND:1 M5:SRC 8.50853e-17 
c_110 GND:1 M17:GATE 9.65559e-19 
c_111 GND:1 M13:GATE 8.38276e-19 
c_112 GND:1 M12:DRN 2.40489e-18 
c_113 GND:1 Q 1.38821e-16 
c_114 GND:1 M4:SRC 2.31157e-18 
c_115 GND:1 E 2.04599e-18 
c_116 GND:1 M7:SRC 1.34823e-18 
c_117 GND:1 M7:GATE 6.22626e-18 
c_118 GND:1 TE 2.37682e-18 
c_119 GND:1 M6:GATE 5.66659e-18 
c_120 GND:1 M5:GATE 4.85928e-18 
c_121 GND:1 0 2.1779e-16 
c_122 M11:SRC Q 5.38077e-18 
c_123 M11:SRC 0 5.45227e-18 
c_124 M14:BULK M5:DRN 8.11588e-18 
c_125 M14:BULK M8:GATE 1.19349e-17 
c_126 M14:BULK M17:GATE 1.19232e-17 
c_127 M14:BULK M18:GATE 9.18063e-18 
c_128 M14:BULK Q 4.86083e-18 
c_129 M14:BULK E 1.69523e-18 
c_130 M14:BULK M7:GATE 1.79835e-17 
c_131 M14:BULK TE 2.99502e-18 
c_132 M14:BULK M6:GATE 5.53123e-18 
c_133 M14:BULK M5:GATE 4.74573e-18 
c_134 M14:BULK M16:DRN 9.45594e-18 
c_135 M14:BULK M27:GATE 8.23549e-18 
c_136 M14:BULK 0 9.07625e-18 
c_137 M14:DRN M5:SRC 2.34847e-22 
c_138 M14:DRN M13:GATE 4.7418e-18 
c_139 M14:DRN M14:SRC 3.97226e-18 
c_140 M14:DRN 0 3.92391e-19 
c_141 M3:DRN M12:DRN 3.05284e-19 
c_142 M3:DRN Q 2.0319e-19 
c_143 M3:DRN 0 9.1122e-18 
c_144 M12:SRC 0 3.91663e-19 
c_145 M4:DRN M4:SRC 3.05284e-19 
c_146 M4:DRN Q 5.57363e-19 
c_147 M4:DRN 0 7.20023e-18 
c_148 M6:SRC M9:SRC 6.59639e-18 
c_149 M6:SRC M5:DRN 1.16348e-17 
c_150 M6:SRC M8:GATE 3.73848e-18 
c_151 M6:SRC M5:SRC 1.44569e-17 
c_152 M6:SRC M17:GATE 5.92967e-19 
c_153 M6:SRC M14:SRC 2.93548e-18 
c_154 M6:SRC M12:DRN 2.92826e-18 
c_155 M6:SRC M4:SRC 2.6162e-18 
c_156 M6:SRC E 2.3443e-19 
c_157 M6:SRC M7:SRC 1.38447e-17 
c_158 M6:SRC M7:GATE 1.85847e-17 
c_159 M6:SRC TE 3.58781e-18 
c_160 M6:SRC M6:GATE 1.80834e-17 
c_161 M6:SRC M5:GATE 8.07105e-18 
c_162 M6:SRC M27:SRC 1.19436e-18 
c_163 M6:SRC M16:DRN 1.78827e-20 
c_164 M6:SRC M1:SRC 1.50098e-18 
c_165 M6:SRC M23:DRN 4.42193e-20 
c_166 M6:SRC M21:DRN 4.42193e-20 
c_167 M6:SRC 0 9.44096e-17 
c_168 GND M7:SRC 1.7848e-20 
c_169 GND E 3.44941e-19 
c_170 GND 0 2.4665e-17 
c_171 M9:DRN M5:DRN 1.78949e-21 
c_172 M9:DRN M8:GATE 2.44177e-17 
c_173 M9:DRN M5:SRC 4.79758e-19 
c_174 M9:DRN M17:GATE 3.11918e-19 
c_175 M9:DRN M15:GATE 1.70314e-19 
c_176 M9:DRN M13:GATE 9.36376e-18 
c_177 M9:DRN M14:SRC 8.09321e-19 
c_178 M9:DRN M12:DRN 3.68254e-19 
c_179 M9:DRN Q 3.34921e-18 
c_180 M9:DRN M4:SRC 3.68254e-19 
c_181 M9:DRN 0 4.37604e-17 
c_182 N_5:1 M9:SRC 1.63588e-18 
c_183 N_5:1 M6:SRC 5.27716e-17 
c_184 N_5:1 M10:GATE 3.90432e-17 
c_185 N_5:1 M19:DRN 3.42234e-19 
c_186 N_5:1 M8:GATE 3.5654e-17 
c_187 N_5:1 M13:DRN 2.1146e-16 
c_188 N_5:1 GND:1 1.73631e-16 
c_189 N_5:1 M9:DRN 9.95117e-18 
c_190 N_5:1 M5:SRC 1.81006e-18 
c_191 N_5:1 M17:GATE 1.18288e-18 
c_192 N_5:1 M18:GATE 3.96596e-17 
c_193 N_5:1 M15:DRN 1.67464e-17 
c_194 N_5:1 M15:GATE 1.67665e-18 
c_195 N_5:1 M13:GATE 4.14952e-18 
c_196 N_5:1 M14:DRN 1.57355e-18 
c_197 N_5:1 M14:BULK 1.51681e-17 
c_198 N_5:1 M14:SRC 6.08747e-17 
c_199 N_5:1 M26:DRN 7.82249e-17 
c_200 N_5:1 M5:GATE 1.19874e-17 
c_201 N_5:1 M1:SRC 4.20333e-18 
c_202 N_5:1 M3:DRN 8.79011e-18 
c_203 N_5:1 0 3.09107e-19 
c_204 M24:GATE GND:1 3.12256e-17 
c_205 M24:GATE M13:GATE 8.53405e-20 
c_206 M24:GATE M16:DRN 5.46435e-21 
c_207 M24:GATE 0 9.85954e-19 
c_208 M1:GATE M6:SRC 1.69314e-18 
c_209 M1:GATE GND:1 5.46035e-18 
c_210 M1:GATE M9:DRN 9.55397e-19 
c_211 M1:GATE M14:BULK 4.59586e-18 
c_212 M1:GATE M3:DRN 1.02864e-17 
c_213 M1:GATE 0 9.97488e-18 
c_214 M18:DRN M6:SRC 6.35686e-20 
c_215 M18:DRN M10:GATE 4.80264e-18 
c_216 M18:DRN M19:DRN 2.12789e-20 
c_217 M18:DRN M8:GATE 2.34862e-18 
c_218 M18:DRN M13:DRN 5.00204e-18 
c_219 M18:DRN GND:1 7.20723e-20 
c_220 M18:DRN M9:DRN 1.01627e-20 
c_221 M18:DRN M17:GATE 3.8456e-18 
c_222 M18:DRN M18:GATE 1.70567e-17 
c_223 M18:DRN M15:DRN 7.41475e-18 
c_224 M18:DRN M15:GATE 6.00903e-18 
c_225 M18:DRN M13:GATE 1.40533e-19 
c_226 M18:DRN M14:BULK 3.44314e-18 
c_227 M18:DRN M14:SRC 2.01118e-20 
c_228 M18:DRN M17:SRC 8.70686e-20 
c_229 M18:DRN M26:DRN 8.00015e-20 
c_230 M18:DRN 0 1.45384e-18 
c_231 M19:GATE M6:SRC 6.45423e-22 
c_232 M19:GATE M8:GATE 7.71572e-18 
c_233 M19:GATE M13:DRN 9.05036e-18 
c_234 M19:GATE M9:DRN 2.41426e-18 
c_235 M19:GATE M17:GATE 9.93101e-18 
c_236 M19:GATE M18:GATE 1.69082e-17 
c_237 M19:GATE M15:DRN 7.10468e-21 
c_238 M19:GATE M15:GATE 4.20697e-21 
c_239 M19:GATE M14:BULK 7.73696e-18 
c_240 M19:GATE M14:SRC 5.51528e-18 
c_241 M19:GATE M17:SRC 2.7673e-18 
c_242 M19:GATE M26:GATE 1.78723e-19 
c_243 M19:GATE M26:DRN 1.63e-19 
c_244 M19:GATE M5:GATE 4.72331e-18 
c_245 M19:GATE 0 9.9795e-19 
c_246 M9:GATE M6:SRC 3.83709e-18 
c_247 M9:GATE M10:GATE 1.02626e-17 
c_248 M9:GATE M8:GATE 1.51546e-17 
c_249 M9:GATE GND:1 4.79516e-18 
c_250 M9:GATE M9:DRN 1.35117e-17 
c_251 M9:GATE M5:SRC 6.50997e-20 
c_252 M9:GATE M14:BULK 4.47892e-18 
c_253 M9:GATE M5:GATE 4.6371e-19 
c_254 M9:GATE 0 1.11012e-17 
c_255 M8:DRN M9:SRC 2.12789e-20 
c_256 M8:DRN M6:SRC 9.42947e-18 
c_257 M8:DRN M8:GATE 1.69748e-17 
c_258 M8:DRN M13:DRN 1.51425e-18 
c_259 M8:DRN GND:1 2.99232e-18 
c_260 M8:DRN M9:DRN 3.41166e-18 
c_261 M8:DRN M5:SRC 8.51908e-20 
c_262 M8:DRN M15:GATE 6.39555e-19 
c_263 M8:DRN M13:GATE 3.932e-18 
c_264 M8:DRN M14:DRN 1.6336e-18 
c_265 M8:DRN M14:SRC 7.80137e-21 
c_266 M8:DRN M12:SRC 3.76568e-22 
c_267 CP:1 M6:SRC 4.5515e-19 
c_268 CP:1 N_5:1 3.29196e-17 
c_269 CP:1 M9:DRN 3.41643e-19 
c_270 CP:1 M13:GATE 3.4497e-17 
c_271 CP:1 M14:BULK 1.74446e-17 
c_272 CP:1 M14:SRC 1.77383e-17 
c_273 CP:1 M1:GATE 7.6789e-18 
c_274 CP:1 M16:DRN 2.3172e-20 
c_275 CP:1 M3:DRN 1.90621e-19 
c_276 CP:1 0 9.44699e-19 
c_277 M25:GATE N_5:1 1.8037e-18 
c_278 M25:GATE M17:GATE 1.17598e-19 
c_279 M25:GATE M15:GATE 2.94769e-19 
c_280 M25:GATE M13:GATE 4.51876e-18 
c_281 M25:GATE M16:DRN 1.70834e-18 
c_282 M25:GATE M24:GATE 8.34247e-18 
c_283 M25:GATE 0 3.00298e-18 
c_284 CP N_5:1 4.62434e-18 
c_285 CP M15:GATE 1.35034e-19 
c_286 CP M13:GATE 1.83474e-17 
c_287 CP M14:BULK 5.83147e-19 
c_288 CP M14:SRC 1.85262e-18 
c_289 CP M16:DRN 7.6603e-17 
c_290 CP 0 4.42303e-18 
c_291 M2:GATE M6:SRC 1.69435e-18 
c_292 M2:GATE N_5:1 6.10898e-18 
c_293 M2:GATE GND:1 1.26932e-18 
c_294 M2:GATE M9:DRN 9.51551e-19 
c_295 M2:GATE M18:DRN 2.78115e-19 
c_296 M2:GATE M13:GATE 1.71123e-19 
c_297 M2:GATE M14:DRN 1.03505e-18 
c_298 M2:GATE M14:BULK 5.61477e-18 
c_299 M2:GATE M14:SRC 1.19401e-19 
c_300 M2:GATE M1:GATE 7.71602e-18 
c_301 M14:GATE M6:SRC 1.99321e-18 
c_302 M14:GATE M8:DRN 7.81739e-20 
c_303 M14:GATE N_5:1 5.39981e-18 
c_304 M14:GATE GND:1 1.19736e-18 
c_305 M14:GATE M9:DRN 7.01386e-19 
c_306 M14:GATE M18:DRN 3.08581e-19 
c_307 M14:GATE M13:GATE 1.01529e-17 
c_308 M14:GATE M14:DRN 1.01125e-17 
c_309 M14:GATE M14:BULK 4.27749e-18 
c_310 M14:GATE M14:SRC 1.52985e-17 
c_311 M14:GATE M1:GATE 5.67619e-20 
c_312 M14:GATE M16:DRN 8.8341e-18 
c_313 M14:GATE 0 5.94781e-18 
c_314 M16:GATE M6:SRC 4.24629e-20 
c_315 M16:GATE N_5:1 5.44382e-19 
c_316 M16:GATE M9:DRN 4.91814e-20 
c_317 M16:GATE M17:GATE 7.53705e-22 
c_318 M16:GATE M18:DRN 1.11446e-18 
c_319 M16:GATE M15:GATE 8.34104e-18 
c_320 M16:GATE M14:DRN 3.06566e-19 
c_321 M16:GATE M16:DRN 2.6694e-17 
c_322 M16:GATE M24:GATE 1.75056e-20 
c_323 M16:GATE 0 8.56139e-18 
c_324 N_13:1 M6:SRC 1.46127e-19 
c_325 N_13:1 N_5:1 1.85245e-16 
c_326 N_13:1 GND:1 3.02829e-18 
c_327 N_13:1 M9:DRN 1.12089e-18 
c_328 N_13:1 M14:BULK 3.14798e-18 
c_329 N_13:1 CP:1 2.8287e-19 
c_330 N_13:1 M1:GATE 1.83575e-17 
c_331 N_13:1 M12:DRN 3.86086e-17 
c_332 N_13:1 Q 5.09811e-17 
c_333 N_13:1 M4:SRC 1.55901e-17 
c_334 N_13:1 M23:DRN 1.44448e-17 
c_335 N_13:1 M21:DRN 1.50154e-17 
c_336 N_13:1 CP 1.56539e-19 
c_337 N_13:1 M25:GATE 1.16914e-19 
c_338 N_13:1 M24:GATE 2.3376e-18 
c_339 N_13:1 M11:SRC 1.72957e-17 
c_340 N_13:1 M3:DRN 6.15561e-18 
c_341 N_13:2 GND:1 6.37163e-18 
c_342 N_13:2 M9:DRN 6.82328e-21 
c_343 N_13:2 M14:BULK 7.99431e-18 
c_344 N_13:2 M1:GATE 8.62901e-20 
c_345 N_13:2 M12:DRN 2.76344e-18 
c_346 N_13:2 Q 1.32513e-17 
c_347 N_13:2 M4:SRC 5.83622e-19 
c_348 N_13:2 M4:DRN 2.62322e-18 
c_349 N_13:2 M24:GATE 6.90321e-20 
c_350 M23:GATE Q 7.75356e-18 
c_351 M23:GATE M23:DRN 3.36346e-17 
c_352 M23:GATE M25:GATE 1.97528e-19 
c_353 M23:GATE M24:GATE 1.05466e-17 
c_354 M23:GATE 0 2.41901e-18 
c_355 M22:GATE Q 2.22486e-17 
c_356 M22:GATE M4:SRC 7.74427e-20 
c_357 M22:GATE M23:DRN 3.34086e-17 
c_358 M22:GATE M21:DRN 2.03258e-19 
c_359 M22:GATE M24:GATE 1.62855e-19 
c_360 M22:GATE 0 5.38129e-19 
c_361 M21:GATE Q 1.70827e-17 
c_362 M21:GATE M23:DRN 2.03258e-19 
c_363 M21:GATE M21:DRN 3.34947e-17 
c_364 M21:GATE 0 2.21354e-18 
c_365 M20:GATE Q 1.07851e-17 
c_366 M20:GATE M4:DRN 3.23339e-18 
c_367 M20:GATE M21:DRN 3.34661e-17 
c_368 M20:GATE 0 1.46566e-18 
c_369 M24:SRC M6:SRC 1.5418e-19 
c_370 M24:SRC N_5:1 2.21136e-17 
c_371 M24:SRC M9:DRN 1.75379e-19 
c_372 M24:SRC M18:DRN 2.35933e-23 
c_373 M24:SRC M15:GATE 3.00857e-17 
c_374 M24:SRC M16:GATE 3.86917e-18 
c_375 M24:SRC M14:BULK 1.52355e-18 
c_376 M24:SRC M14:SRC 5.4886e-19 
c_377 M24:SRC CP:1 9.01582e-18 
c_378 M24:SRC M2:GATE 4.26731e-18 
c_379 M24:SRC M16:DRN 7.98401e-19 
c_380 M24:SRC M1:SRC 4.62556e-19 
c_381 M24:SRC M23:DRN 4.05118e-20 
c_382 M24:SRC CP 8.23601e-17 
c_383 M24:SRC M25:GATE 2.90092e-17 
c_384 M24:SRC M24:GATE 1.84318e-17 
c_385 M24:SRC 0 3.2797e-19 
c_386 M4:GATE M6:SRC 1.73264e-18 
c_387 M4:GATE GND:1 7.72197e-18 
c_388 M4:GATE M9:DRN 1.09704e-18 
c_389 M4:GATE M14:BULK 6.34968e-18 
c_390 M4:GATE M12:SRC 1.84847e-18 
c_391 M4:GATE Q 3.34185e-18 
c_392 M4:GATE M4:SRC 1.67248e-17 
c_393 M4:GATE M4:DRN 1.08873e-17 
c_394 M11:GATE M4:SRC 1.60344e-17 
c_395 M11:GATE Q 9.56804e-19 
c_396 M11:GATE GND:1 4.14686e-18 
c_397 M11:GATE M14:BULK 3.3432e-18 
c_398 M11:GATE M12:DRN 7.74427e-20 
c_399 M11:GATE M12:SRC 8.3794e-18 
c_400 M11:GATE M6:SRC 1.74486e-18 
c_401 M11:GATE M9:DRN 8.66301e-18 
c_402 M12:GATE M6:SRC 2.04938e-18 
c_403 M12:GATE GND:1 5.21656e-18 
c_404 M12:GATE M9:DRN 8.4051e-18 
c_405 M12:GATE M14:BULK 4.03502e-18 
c_406 M12:GATE M1:GATE 8.83887e-20 
c_407 M12:GATE M12:DRN 7.4765e-18 
c_408 M12:GATE M12:SRC 8.33984e-18 
c_409 M12:GATE Q 1.06756e-17 
c_410 M12:GATE M3:DRN 1.2593e-20 
c_411 M3:GATE M6:SRC 1.73264e-18 
c_412 M3:GATE N_5:1 3.42457e-20 
c_413 M3:GATE GND:1 7.97358e-18 
c_414 M3:GATE M9:DRN 1.09704e-18 
c_415 M3:GATE M14:BULK 3.96449e-18 
c_416 M3:GATE CP:1 9.16955e-21 
c_417 M3:GATE M2:GATE 4.81174e-19 
c_418 M3:GATE M1:GATE 5.92707e-18 
c_419 M3:GATE M12:SRC 1.84847e-18 
c_420 M3:GATE Q 1.28635e-18 
c_421 M3:GATE M24:GATE 7.41991e-19 
c_422 M3:GATE M3:DRN 1.66894e-17 
c_423 M3:GATE 0 1.47119e-18 
c_424 M2:SRC M6:SRC 2.84478e-18 
c_425 M2:SRC N_5:1 3.86816e-18 
c_426 M2:SRC GND:1 2.36512e-17 
c_427 M2:SRC M9:DRN 4.53683e-19 
c_428 M2:SRC M13:GATE 1.1805e-18 
c_429 M2:SRC M14:DRN 2.17028e-20 
c_430 M2:SRC M14:SRC 2.02535e-17 
c_431 M2:SRC CP:1 2.06842e-17 
c_432 M2:SRC M2:GATE 1.44945e-17 
c_433 M2:SRC M1:GATE 1.22902e-18 
c_434 M2:SRC M12:DRN 4.63261e-19 
c_435 M2:SRC Q 8.55661e-17 
c_436 M2:SRC M23:DRN 1.20032e-18 
c_437 M2:SRC CP 8.1805e-19 
c_438 M2:SRC M24:GATE 6.19557e-18 
c_439 M2:SRC M3:DRN 1.62168e-18 
c_440 M2:SRC 0 1.39569e-17 
c_441 VDD:1 N_5:1 2.99625e-19 
c_442 VDD:1 M17:GATE 1.15837e-18 
c_443 VDD:1 M19:GATE 5.06722e-19 
c_444 VDD:1 M18:GATE 1.94689e-20 
c_445 VDD:1 M15:DRN 4.29761e-19 
c_446 VDD:1 M15:GATE 7.90313e-18 
c_447 VDD:1 M16:GATE 5.69847e-18 
c_448 VDD:1 M14:GATE 7.13088e-19 
c_449 VDD:1 M24:SRC 6.77174e-18 
c_450 VDD:1 Q 1.24699e-17 
c_451 VDD:1 M26:GATE 3.6792e-17 
c_452 VDD:1 M16:DRN 5.88873e-17 
c_453 VDD:1 M27:GATE 1.15091e-19 
c_454 VDD:1 CP 3.37452e-18 
c_455 VDD:1 M25:GATE 2.47445e-18 
c_456 VDD:1 M24:GATE 6.53728e-19 
c_457 VDD:1 M22:GATE 7.63052e-19 
c_458 VDD:1 M23:GATE 1.28696e-18 
c_459 VDD:1 0 3.56919e-17 
c_460 VDD:2 N_5:1 3.78688e-19 
c_461 VDD:2 M17:GATE 2.89828e-19 
c_462 VDD:2 M13:GATE 7.38557e-19 
c_463 VDD:2 M16:GATE 8.35541e-20 
c_464 VDD:2 M2:SRC 3.21953e-17 
c_465 VDD:2 M24:SRC 3.98679e-19 
c_466 VDD:2 N_13:1 1.13755e-18 
c_467 VDD:2 Q 9.73399e-17 
c_468 VDD:2 M23:DRN 1.53596e-19 
c_469 VDD:2 M21:DRN 7.33167e-19 
c_470 VDD:2 M25:GATE 1.96167e-18 
c_471 VDD:2 M24:GATE 4.00231e-18 
c_472 VDD:2 M20:GATE 9.26983e-18 
c_473 VDD:2 M22:GATE 1.72859e-18 
c_474 VDD:2 M21:GATE 3.08658e-18 
c_475 VDD:2 M23:GATE 1.44255e-18 
c_476 VDD:2 0 2.78076e-17 
c_477 M25:BULK M10:GATE 1.35083e-17 
c_478 M25:BULK M8:GATE 9.12926e-19 
c_479 M25:BULK N_5:1 1.11224e-17 
c_480 M25:BULK M13:DRN 1.13648e-17 
c_481 M25:BULK M17:GATE 2.11854e-17 
c_482 M25:BULK M19:GATE 4.41373e-19 
c_483 M25:BULK M9:GATE 3.682e-18 
c_484 M25:BULK M18:GATE 6.15153e-18 
c_485 M25:BULK M18:DRN 2.51369e-18 
c_486 M25:BULK M15:DRN 1.6422e-18 
c_487 M25:BULK M15:GATE 1.09983e-17 
c_488 M25:BULK M13:GATE 9.61703e-18 
c_489 M25:BULK M16:GATE 1.40519e-17 
c_490 M25:BULK M14:SRC 2.97489e-25 
c_491 M25:BULK CP:1 6.50026e-19 
c_492 M25:BULK M24:SRC 7.38926e-18 
c_493 M25:BULK N_13:1 2.08254e-19 
c_494 M25:BULK Q 6.41023e-18 
c_495 M25:BULK N_13:2 8.56215e-18 
c_496 M25:BULK E 6.55934e-18 
c_497 M25:BULK TE 5.06942e-18 
c_498 M25:BULK M6:GATE 3.59496e-18 
c_499 M25:BULK M26:GATE 4.54509e-18 
c_500 M25:BULK M26:DRN 3.08152e-18 
c_501 M25:BULK M23:DRN 3.656e-18 
c_502 M25:BULK M21:DRN 2.40244e-18 
c_503 M25:BULK M27:GATE 5.09848e-18 
c_504 M25:BULK M25:GATE 1.32633e-17 
c_505 M25:BULK M24:GATE 2.98019e-18 
c_506 M25:BULK M28:GATE 1.01211e-17 
c_507 M25:BULK M20:GATE 7.23515e-18 
c_508 M25:BULK M22:GATE 3.55168e-18 
c_509 M25:BULK M21:GATE 3.87465e-18 
c_510 M25:BULK M23:GATE 4.77326e-18 
c_511 VDD M10:GATE 5.18663e-17 
c_512 VDD N_5:1 3.11584e-18 
c_513 VDD M5:SRC 2.00372e-18 
c_514 VDD M17:GATE 4.38696e-17 
c_515 VDD M18:GATE 1.25481e-18 
c_516 VDD M18:DRN 8.30063e-19 
c_517 VDD M15:DRN 1.20574e-16 
c_518 VDD M15:GATE 1.85601e-18 
c_519 VDD M16:GATE 1.34043e-18 
c_520 VDD M14:SRC 1.2687e-17 
c_521 VDD CP:1 1.42513e-20 
c_522 VDD M24:SRC 1.88822e-18 
c_523 VDD N_13:1 1.59292e-17 
c_524 VDD Q 4.29773e-17 
c_525 VDD E 3.52891e-17 
c_526 VDD TE 2.68863e-17 
c_527 VDD M26:GATE 6.08601e-18 
c_528 VDD M26:DRN 1.34853e-18 
c_529 VDD M27:SRC 5.10732e-19 
c_530 VDD M26:SRC 3.62831e-19 
c_531 VDD M16:DRN 1.59769e-18 
c_532 VDD M23:DRN 2.66033e-18 
c_533 VDD M21:DRN 2.66033e-18 
c_534 VDD M27:GATE 8.71193e-18 
c_535 VDD CP 1.61747e-19 
c_536 VDD M25:GATE 5.22944e-18 
c_537 VDD M24:GATE 4.39694e-18 
c_538 VDD M28:GATE 1.33601e-17 
c_539 VDD M20:GATE 3.71611e-18 
c_540 VDD M22:GATE 3.79346e-18 
c_541 VDD M21:GATE 4.47108e-18 
c_542 VDD M23:GATE 4.61683e-18 
c_543 VDD 0 1.83264e-16 
c_544 M16:SRC M10:GATE 2.75143e-18 
c_545 M16:SRC M8:GATE 6.10875e-19 
c_546 M16:SRC M8:DRN 1.0157e-19 
c_547 M16:SRC N_5:1 4.03594e-19 
c_548 M16:SRC M13:DRN 5.91887e-20 
c_549 M16:SRC M5:SRC 1.08052e-19 
c_550 M16:SRC M17:GATE 1.09454e-16 
c_551 M16:SRC M19:GATE 2.39037e-19 
c_552 M16:SRC M18:GATE 7.79826e-19 
c_553 M16:SRC M18:DRN 9.81936e-19 
c_554 M16:SRC M15:DRN 9.56395e-18 
c_555 M16:SRC M15:GATE 5.38379e-17 
c_556 M16:SRC M16:GATE 2.77088e-17 
c_557 M16:SRC M14:SRC 7.22355e-18 
c_558 M16:SRC M2:SRC 7.81718e-21 
c_559 M16:SRC CP:1 1.28377e-19 
c_560 M16:SRC M24:SRC 8.85823e-18 
c_561 M16:SRC N_13:1 6.58196e-20 
c_562 M16:SRC M12:DRN 3.81007e-20 
c_563 M16:SRC M4:SRC 3.81007e-20 
c_564 M16:SRC M17:SRC 7.4898e-18 
c_565 M16:SRC E 1.01891e-19 
c_566 M16:SRC TE 7.3625e-19 
c_567 M16:SRC M26:GATE 9.50019e-18 
c_568 M16:SRC M26:DRN 1.08701e-18 
c_569 M16:SRC M27:SRC 6.53413e-18 
c_570 M16:SRC M26:SRC 6.52944e-18 
c_571 M16:SRC M16:DRN 1.13799e-17 
c_572 M16:SRC M23:DRN 1.00992e-17 
c_573 M16:SRC M21:DRN 1.00992e-17 
c_574 M16:SRC M27:GATE 9.5041e-18 
c_575 M16:SRC M25:GATE 4.88646e-18 
c_576 M16:SRC M24:GATE 4.35799e-18 
c_577 M16:SRC M28:GATE 9.50033e-18 
c_578 M16:SRC M20:GATE 4.35799e-18 
c_579 M16:SRC M22:GATE 5.29123e-18 
c_580 M16:SRC M21:GATE 4.35799e-18 
c_581 M16:SRC M23:GATE 4.35799e-18 
c_582 M16:SRC 0 1.34366e-16 
c_583 M22:DRN Q 1.90512e-17 
c_584 M22:DRN N_13:1 1.4812e-17 
c_585 M22:DRN M23:GATE 9.20638e-19 
c_586 M22:DRN M22:GATE 2.09805e-17 
c_587 M22:DRN M21:GATE 2.06656e-17 
c_588 M22:DRN M20:GATE 1.97061e-18 
c_589 M22:DRN 0 5.92181e-18 
c_590 M25:SRC N_5:1 3.46254e-20 
c_591 M25:SRC M17:GATE 8.61901e-19 
c_592 M25:SRC M18:DRN 3.37527e-21 
c_593 M25:SRC M15:GATE 4.42618e-19 
c_594 M25:SRC M13:GATE 8.1852e-19 
c_595 M25:SRC M16:GATE 5.1165e-18 
c_596 M25:SRC M14:GATE 4.40112e-18 
c_597 M25:SRC M2:SRC 4.20236e-19 
c_598 M25:SRC CP:1 9.87393e-21 
c_599 M25:SRC M24:SRC 1.50085e-18 
c_600 M25:SRC N_13:1 1.00965e-19 
c_601 M25:SRC Q 1.74812e-18 
c_602 M25:SRC M26:GATE 6.04706e-20 
c_603 M25:SRC M16:DRN 1.7902e-17 
c_604 M25:SRC M23:DRN 8.45673e-19 
c_605 M25:SRC M21:DRN 8.45673e-19 
c_606 M25:SRC CP 3.86637e-19 
c_607 M25:SRC M25:GATE 2.49372e-17 
c_608 M25:SRC M24:GATE 6.69023e-18 
c_609 M25:SRC M20:GATE 5.14009e-18 
c_610 M25:SRC M22:GATE 3.76889e-18 
c_611 M25:SRC M21:GATE 5.1394e-18 
c_612 M25:SRC M23:GATE 5.14089e-18 
c_613 M25:SRC 0 1.55411e-17 
c_614 M24:DRN M2:SRC 6.38043e-18 
c_615 M24:DRN N_13:1 1.05663e-19 
c_616 M24:DRN Q 2.36314e-19 
c_617 M24:DRN M23:DRN 4.61361e-19 
c_618 M24:DRN M25:GATE 9.39271e-19 
c_619 M24:DRN M24:GATE 2.76274e-17 
c_620 M24:DRN M22:GATE 1.44143e-18 
c_621 M24:DRN M23:GATE 2.87138e-17 
c_622 M24:DRN 0 5.71548e-19 
c_623 M23:SRC N_13:1 5.11979e-18 
c_624 M23:SRC N_5:1 9.78277e-18 
c_625 M23:SRC M25:GATE 1.32985e-18 
c_626 M23:SRC M24:GATE 5.71774e-18 
c_627 M23:SRC M2:SRC 2.36229e-18 
c_628 M23:SRC M18:DRN 1.28891e-19 
c_629 M23:SRC 0 5.50281e-18 
c_630 M20:DRN M20:GATE 3.51846e-17 
c_631 M20:DRN M21:DRN 1.50316e-18 
c_632 M20:DRN M21:GATE 4.4775e-20 
c_633 M20:DRN Q 1.11495e-18 
c_634 M20:DRN 0 6.27607e-18 
c_635 M28:SRC M26:SRC 6.57189e-19 
c_636 M28:SRC M27:GATE 3.21378e-19 
c_637 M28:SRC M28:GATE 3.39622e-17 
c_638 M28:SRC E 2.1928e-17 
c_639 M28:SRC TE 1.1937e-19 
c_640 M28:SRC 0 8.99865e-19 
c_641 M19:SRC M10:GATE 5.8544e-18 
c_642 M19:SRC N_5:1 1.62116e-18 
c_643 M19:SRC M17:GATE 9.06424e-18 
c_644 M19:SRC M19:GATE 1.99137e-17 
c_645 M19:SRC M18:GATE 7.88108e-18 
c_646 M19:SRC M15:DRN 1.87971e-18 
c_647 M19:SRC M15:GATE 2.85073e-17 
c_648 M19:SRC M16:GATE 4.38482e-21 
c_649 M19:SRC M17:SRC 1.32064e-17 
c_650 M19:SRC M26:GATE 2.79519e-19 
c_651 M19:SRC M5:GATE 7.12028e-19 
c_652 M19:SRC M26:SRC 2.22238e-20 
c_653 M19:SRC 0 2.51125e-18 

.ENDS
