
.subckt CKBD8  CLK C
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.07452p as=0.05589p l=0.09u nrd=0.572 nrs=0.431 pd=0.891u ps=0.6642u sa=6.21e-07 sb=2.502e-06 w=0.36u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.04212p as=0.08181p l=0.09u nrd=0.325 nrs=0.629 pd=0.594u ps=0.882u sa=2.52e-06 sb=6.03e-07 w=0.36u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.04212p as=0.08181p l=0.09u nrd=0.325 nrs=0.629 pd=0.594u ps=0.882u sa=1.782e-06 sb=1.341e-06 w=0.36u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.04212p as=0.07452p l=0.09u nrd=0.325 nrs=0.572 pd=0.594u ps=0.891u sa=1.044e-06 sb=2.079e-06 w=0.36u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.13365p as=0.06966p l=0.09u nrd=0.661 nrs=0.344 pd=1.764u ps=0.8298u sa=2.34e-07 sb=8.928e-07 w=0.45u 
DDD1 DD1:ANODE DD1:CATHODE ndio area=0.081p pj=1.26u
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.14661p as=0.04212p l=0.09u nrd=1.133 nrs=0.325 pd=1.674u ps=0.594u sa=2.844e-06 sb=2.79e-07 w=0.36u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.08181p as=0.04212p l=0.09u nrd=0.629 nrs=0.325 pd=0.882u ps=0.594u sa=2.106e-06 sb=1.017e-06 w=0.36u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.08181p as=0.04212p l=0.09u nrd=0.629 nrs=0.325 pd=0.882u ps=0.594u sa=1.368e-06 sb=1.755e-06 w=0.36u 
MM9 M9:DRN M9:GATE M9:SRC M9:BULK pch ad=0.08424p as=0.08262p l=0.09u nrd=0.65 nrs=0.637 pd=1.188u ps=0.8127u sa=3.528e-06 sb=2.34e-07 w=0.36u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK pch ad=0.20655p as=0.1053p l=0.09u nrd=0.255 nrs=0.13 pd=2.0313u ps=1.134u sa=2.7666e-06 sb=3.168e-07 w=0.9u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK pch ad=0.14418p as=0.1053p l=0.09u nrd=0.178 nrs=0.13 pd=1.377u ps=1.134u sa=2.025e-06 sb=1.0575e-06 w=0.9u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK pch ad=0.13932p as=0.1053p l=0.09u nrd=0.172 nrs=0.13 pd=1.368u ps=1.134u sa=1.2114e-06 sb=1.7541e-06 w=0.9u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK pch ad=0.14742p as=0.08424p l=0.09u nrd=0.284 nrs=0.162 pd=1.3041u ps=0.954u sa=9.54e-07 sb=2.592e-06 w=0.72u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK pch ad=0.16848p as=0.12474p l=0.09u nrd=0.325 nrs=0.24 pd=1.908u ps=1.224u sa=2.34e-07 sb=3.3147e-06 w=0.72u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK pch ad=0.1053p as=0.14418p l=0.09u nrd=0.13 nrs=0.178 pd=1.134u ps=1.377u sa=2.4246e-06 sb=6.732e-07 w=0.9u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK pch ad=0.1053p as=0.13932p l=0.09u nrd=0.13 nrs=0.172 pd=1.134u ps=1.368u sa=1.6578e-06 sb=1.3887e-06 w=0.9u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK pch ad=0.1053p as=0.18387p l=0.09u nrd=0.13 nrs=0.227 pd=1.134u ps=1.6299u sa=7.002e-07 sb=2.0817e-06 w=0.9u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK pch ad=0.08424p as=0.12474p l=0.09u nrd=0.162 nrs=0.24 pd=0.954u ps=1.224u sa=6.3e-07 sb=2.9178e-06 w=0.72u 
R1 CLK:1 M8:GATE 58.92
R2 CLK:1 M7:GATE 86.6992
R3 CLK:1 M16:GATE 93.8163
R4 CLK:1 CLK 37.4388
R5 CLK:1 M18:GATE 120.379
R6 CLK:1 M17:GATE 69.6
R7 M18:GATE CLK 216.313
R8 M16:GATE M7:GATE 518.819
R9 CLK DD1:CATHODE 18.1388
R10 GND:1 M4:SRC 18
R11 GND:1 M6:SRC 18.6298
R12 GND:1 M8:DRN 1.28509
R13 GND:1 GND 0.32049
R14 GND M8:DRN 3.7353
R15 M2:SRC M3:DRN 0.001
R16 M2:SRC M8:DRN 2.38411e-10
R17 M8:DRN M4:SRC 0.001
R18 M8:DRN M6:SRC 0.001
R19 M8:DRN DD1:ANODE 0.001
R20 M8:DRN M8:BULK 0.001
R21 M8:DRN M7:BULK 0.001
R22 M8:DRN M6:BULK 0.001
R23 M8:DRN M5:BULK 0.001
R24 M8:DRN M4:BULK 0.001
R25 M8:DRN M3:BULK 0.001
R26 M8:DRN M2:BULK 0.001
R27 M8:DRN M1:BULK 0.001
R28 M8:DRN M1:DRN 0.001
R29 M6:SRC M7:DRN 0.001
R30 M4:SRC M5:DRN 0.001
R31 C:1 C 0.285829
R32 C:1 M15:DRN 23.4593
R33 C:1 M13:DRN 23.4296
R34 C:1 M11:DRN 9.00001
R35 C:1 M9:DRN 18.3458
R36 M11:DRN M10:SRC 0.001
R37 C M4:DRN 18.2456
R38 C M5:SRC 18.4902
R39 C M1:SRC 18.5351
R40 C M15:DRN 15.2716
R41 C M13:DRN 14.9665
R42 M1:SRC M2:DRN 0.001
R43 M4:DRN M3:SRC 0.001
R44 M15:DRN M14:SRC 0.001
R45 M13:DRN M12:SRC 0.001
R46 M5:SRC M6:DRN 0.001
R47 N_12:1 N_12:2 18.0462
R48 N_12:1 M2:GATE 45.36
R49 N_12:1 M1:GATE 79.5618
R50 N_12:1 M11:GATE 77.76
R51 N_12:1 M10:GATE 136.392
R52 N_12:1 M9:GATE 187.247
R53 N_12:2 N_12:5 42.3665
R54 N_12:2 M4:GATE 104.564
R55 N_12:2 M3:GATE 31.32
R56 N_12:2 M13:GATE 181.415
R57 N_12:2 M12:GATE 63.72
R58 N_12:3 N_12:5 13.4334
R59 N_12:3 N_12:4 16.4277
R60 N_12:3 M7:SRC 1175.61
R61 N_12:3 M6:GATE 33.0109
R62 N_12:3 M15:GATE 72.2109
R63 N_12:4 N_12:5 16.5945
R64 N_12:4 M7:SRC 18.9994
R65 N_12:4 M18:DRN 9.60983
R66 N_12:4 M17:DRN 9.13048
R67 M10:GATE M1:GATE 363.268
R68 M10:GATE M9:GATE 854.943
R69 M9:GATE M1:GATE 498.717
R70 N_12:5 M7:SRC 1187.54
R71 N_12:5 M5:GATE 33.5082
R72 N_12:5 M4:GATE 124.896
R73 N_12:5 M14:GATE 72.7082
R74 N_12:5 M13:GATE 216.69
R75 M4:GATE M13:GATE 534.807
R76 M17:DRN M16:SRC 0.001
R77 M7:SRC M8:SRC 0.001
R78 VDD:1 M18:SRC 2.6009
R79 VDD:1 M14:DRN 18
R80 VDD:1 M16:DRN 14.966
R81 VDD:1 VDD 0.324226
R82 VDD:1 VDD:2 0.237777
R83 VDD:2 M18:SRC 3.49158
R84 VDD:2 M12:DRN 18.3054
R85 VDD:2 M10:DRN 18
R86 VDD M18:SRC 3.18386
R87 VDD M16:DRN 25.8976
R88 M12:DRN M18:SRC 9.52381e-11
R89 M12:DRN M11:SRC 0.001
R90 M10:DRN M18:SRC 7.69231e-11
R91 M10:DRN M9:SRC 0.001
R92 M14:DRN M18:SRC 4.08064e-10
R93 M14:DRN M13:SRC 0.001
R94 M18:SRC M16:DRN 4.9537e-10
R95 M18:SRC M17:SRC 0.001
R96 M18:SRC M18:BULK 0.001
R97 M18:SRC M17:BULK 0.001
R98 M18:SRC M16:BULK 0.001
R99 M18:SRC M15:BULK 0.001
R100 M18:SRC M14:BULK 0.001
R101 M18:SRC M13:BULK 0.001
R102 M18:SRC M12:BULK 0.001
R103 M18:SRC M11:BULK 0.001
R104 M18:SRC M10:BULK 0.001
R105 M18:SRC M9:BULK 0.001
R106 M16:DRN M15:SRC 0.001
c_1 CLK:1 0 5.29485e-19 
c_2 M18:GATE 0 2.77076e-17 
c_3 M17:GATE 0 1.07841e-18 
c_4 M16:GATE 0 9.1312e-19 
c_5 CLK 0 7.98451e-18 
c_6 M8:GATE 0 7.29415e-21 
c_7 M7:GATE 0 1.713e-19 
c_8 DD1:CATHODE 0 9.37659e-19 
c_9 GND:1 CLK:1 4.2457e-18 
c_10 GND:1 M8:GATE 1.02281e-17 
c_11 GND:1 M7:GATE 8.85522e-18 
c_12 GND:1 CLK 1.69756e-17 
c_13 GND:1 DD1:CATHODE 1.62472e-18 
c_14 GND:1 0 1.69694e-16 
c_15 GND CLK:1 3.30595e-21 
c_16 GND CLK 1.83605e-17 
c_17 GND M7:GATE 5.14814e-19 
c_18 GND DD1:CATHODE 8.17113e-21 
c_19 GND 0 5.042e-17 
c_20 M2:SRC 0 5.72551e-18 
c_21 M8:DRN CLK:1 4.78056e-17 
c_22 M8:DRN M8:GATE 2.40044e-17 
c_23 M8:DRN M7:GATE 1.34178e-17 
c_24 M8:DRN CLK 1.06296e-17 
c_25 M8:DRN DD1:CATHODE 2.82226e-17 
c_26 M8:DRN 0 8.96257e-17 
c_27 M6:SRC CLK:1 1.04135e-18 
c_28 M6:SRC M8:GATE 1.16401e-18 
c_29 M6:SRC M7:GATE 1.19906e-17 
c_30 M6:SRC M16:GATE 8.03616e-18 
c_31 M6:SRC 0 1.10235e-17 
c_32 M4:SRC 0 1.17382e-17 
c_33 C:1 0 4.62239e-17 
c_34 C M4:SRC 7.86034e-18 
c_35 C M6:SRC 4.30058e-19 
c_36 C M8:DRN 5.52236e-17 
c_37 C GND:1 1.48058e-16 
c_38 C GND 2.27301e-17 
c_39 C M2:SRC 5.93853e-18 
c_40 C 0 8.5055e-19 
c_41 M9:DRN GND:1 1.66351e-18 
c_42 M9:DRN M8:DRN 2.03015e-18 
c_43 M9:DRN 0 5.26007e-19 
c_44 M1:SRC M8:DRN 1.00908e-17 
c_45 M1:SRC GND:1 2.55171e-18 
c_46 M1:SRC 0 1.73959e-18 
c_47 M4:DRN M8:DRN 9.11855e-18 
c_48 M4:DRN GND:1 2.24158e-18 
c_49 M4:DRN 0 1.66983e-18 
c_50 M15:DRN M8:DRN 4.17822e-21 
c_51 M15:DRN 0 6.56324e-18 
c_52 M13:DRN 0 2.4491e-18 
c_53 M5:SRC M6:SRC 2.03163e-19 
c_54 M5:SRC M8:DRN 1.05906e-17 
c_55 M5:SRC GND:1 2.64726e-18 
c_56 M5:SRC 0 1.75614e-18 
c_57 N_12:1 M8:DRN 6.38451e-18 
c_58 N_12:1 GND:1 1.44354e-18 
c_59 N_12:1 C 8.4918e-18 
c_60 N_12:1 M1:SRC 1.45577e-17 
c_61 N_12:1 M13:DRN 1.44835e-19 
c_62 N_12:1 M11:DRN 5.93478e-17 
c_63 N_12:1 C:1 1.38517e-17 
c_64 N_12:2 M4:DRN 3.34329e-17 
c_65 N_12:2 M4:SRC 2.2207e-17 
c_66 N_12:2 M5:SRC 1.66747e-17 
c_67 N_12:2 M8:DRN 3.84402e-17 
c_68 N_12:2 CLK:1 1.92055e-18 
c_69 N_12:2 GND:1 1.0887e-17 
c_70 N_12:2 C 8.42491e-17 
c_71 N_12:2 M1:SRC 1.63755e-17 
c_72 N_12:2 M8:GATE 1.10078e-20 
c_73 N_12:2 M7:GATE 3.29303e-18 
c_74 N_12:2 CLK 2.84063e-20 
c_75 N_12:2 M15:DRN 1.97867e-17 
c_76 N_12:2 M13:DRN 1.83045e-17 
c_77 N_12:2 M2:SRC 2.05914e-17 
c_78 N_12:2 M11:DRN 1.96624e-17 
c_79 N_12:3 M4:SRC 1.90572e-20 
c_80 N_12:3 M5:SRC 5.38946e-18 
c_81 N_12:3 M6:SRC 8.78705e-18 
c_82 N_12:3 M8:DRN 1.51805e-18 
c_83 N_12:3 CLK:1 1.54417e-18 
c_84 N_12:3 GND:1 5.41384e-19 
c_85 N_12:3 C 4.6767e-18 
c_86 N_12:3 M8:GATE 9.28231e-20 
c_87 N_12:3 M7:GATE 1.0656e-18 
c_88 N_12:3 M16:GATE 1.20975e-18 
c_89 N_12:3 CLK 3.66383e-20 
c_90 N_12:3 GND 3.45248e-18 
c_91 N_12:3 0 4.37877e-18 
c_92 N_12:4 M4:SRC 4.45877e-19 
c_93 N_12:4 M5:SRC 1.13985e-18 
c_94 N_12:4 M6:SRC 3.07194e-18 
c_95 N_12:4 M8:DRN 3.35983e-17 
c_96 N_12:4 CLK:1 2.1627e-17 
c_97 N_12:4 GND:1 8.99561e-17 
c_98 N_12:4 C 9.22368e-17 
c_99 N_12:4 M8:GATE 4.86333e-18 
c_100 N_12:4 M7:GATE 4.10626e-18 
c_101 N_12:4 M16:GATE 1.50669e-19 
c_102 N_12:4 CLK 9.85245e-17 
c_103 N_12:4 DD1:CATHODE 3.87864e-19 
c_104 N_12:4 GND 2.49076e-19 
c_105 N_12:4 M15:DRN 1.06512e-18 
c_106 N_12:4 M13:DRN 1.38722e-20 
c_107 N_12:4 M11:DRN 1.38722e-20 
c_108 N_12:4 M18:GATE 1.49891e-19 
c_109 N_12:4 C:1 1.43801e-18 
c_110 N_12:4 M17:GATE 1.01962e-17 
c_111 N_12:4 0 1.71699e-17 
c_112 M11:GATE C:1 7.78806e-18 
c_113 M11:GATE M11:DRN 1.042e-17 
c_114 M10:GATE M1:SRC 1.37991e-17 
c_115 M10:GATE M11:DRN 1.27931e-18 
c_116 M10:GATE M9:DRN 2.23067e-19 
c_117 M10:GATE C:1 3.34531e-18 
c_118 M10:GATE 0 3.55922e-18 
c_119 M9:GATE C:1 1.036e-17 
c_120 M9:GATE M11:DRN 3.94166e-19 
c_121 M9:GATE M9:DRN 1.65576e-17 
c_122 M9:GATE 0 8.68627e-18 
c_123 N_12:5 M4:DRN 9.47617e-18 
c_124 N_12:5 M4:SRC 6.12473e-22 
c_125 N_12:5 M5:SRC 1.05606e-17 
c_126 N_12:5 M6:SRC 1.34276e-20 
c_127 N_12:5 M8:DRN 1.96866e-18 
c_128 N_12:5 CLK:1 7.23146e-20 
c_129 N_12:5 GND:1 1.29436e-18 
c_130 N_12:5 C 1.24549e-17 
c_131 N_12:5 M15:DRN 2.07391e-21 
c_132 M4:GATE C 8.47164e-18 
c_133 M4:GATE GND:1 4.8834e-18 
c_134 M4:GATE M4:DRN 3.60111e-18 
c_135 M4:GATE M8:DRN 1.49077e-17 
c_136 M4:GATE M4:SRC 1.78321e-17 
c_137 M4:GATE M5:SRC 4.97775e-20 
c_138 M4:GATE 0 1.99732e-18 
c_139 M2:GATE GND:1 5.01039e-18 
c_140 M2:GATE C 8.3245e-18 
c_141 M2:GATE M1:SRC 3.21277e-18 
c_142 M2:GATE M4:DRN 1.08817e-19 
c_143 M2:GATE M8:DRN 3.26477e-17 
c_144 M1:GATE GND:1 8.54567e-18 
c_145 M1:GATE C 1.54189e-19 
c_146 M1:GATE C:1 1.46735e-17 
c_147 M1:GATE M1:SRC 2.96369e-18 
c_148 M1:GATE M8:DRN 4.39877e-17 
c_149 M15:GATE CLK:1 1.03991e-18 
c_150 M15:GATE C 8.16356e-18 
c_151 M15:GATE M16:GATE 3.89864e-18 
c_152 M15:GATE CLK 8.17961e-20 
c_153 M15:GATE M15:DRN 3.29105e-17 
c_154 M15:GATE C:1 2.40735e-18 
c_155 M15:GATE M17:GATE 1.8914e-19 
c_156 M15:GATE 0 1.37349e-18 
c_157 M14:GATE CLK:1 7.11998e-20 
c_158 M14:GATE C 9.21106e-18 
c_159 M14:GATE M16:GATE 1.64415e-19 
c_160 M14:GATE M15:DRN 3.44553e-17 
c_161 M14:GATE M13:DRN 1.54885e-19 
c_162 M14:GATE C:1 8.12124e-18 
c_163 M14:GATE 0 2.49311e-19 
c_164 M13:GATE C 1.74101e-20 
c_165 M13:GATE M15:DRN 1.54885e-19 
c_166 M13:GATE M13:DRN 3.44753e-17 
c_167 M13:GATE C:1 2.36524e-17 
c_168 M13:GATE 0 1.82852e-18 
c_169 M12:GATE M13:DRN 3.43728e-17 
c_170 M12:GATE M11:DRN 1.44835e-19 
c_171 M12:GATE C:1 2.6404e-17 
c_172 M12:GATE 0 4.71333e-19 
c_173 M18:DRN CLK:1 4.73198e-17 
c_174 M18:DRN CLK 1.17561e-18 
c_175 M18:DRN DD1:CATHODE 2.27425e-18 
c_176 M18:DRN 0 1.07745e-17 
c_177 M17:DRN CLK:1 5.23583e-17 
c_178 M17:DRN CLK 1.5059e-17 
c_179 M17:DRN M15:DRN 5.71598e-20 
c_180 M17:DRN M17:GATE 1.61973e-17 
c_181 M17:DRN 0 2.06831e-18 
c_182 M5:GATE C 4.58327e-19 
c_183 M5:GATE M4:DRN 1.08817e-19 
c_184 M5:GATE GND:1 4.91738e-18 
c_185 M5:GATE M7:GATE 1.44992e-19 
c_186 M5:GATE M8:DRN 1.25446e-17 
c_187 M5:GATE M6:SRC 1.16158e-18 
c_188 M5:GATE M4:SRC 1.8158e-17 
c_189 M5:GATE M5:SRC 6.15431e-18 
c_190 M6:GATE C 1.54318e-19 
c_191 M6:GATE GND:1 4.71422e-18 
c_192 M6:GATE M7:GATE 1.14825e-18 
c_193 M6:GATE M8:GATE 1.39784e-19 
c_194 M6:GATE M8:DRN 1.2647e-17 
c_195 M6:GATE M6:SRC 9.64992e-18 
c_196 M6:GATE M4:SRC 1.19815e-18 
c_197 M6:GATE M5:SRC 1.1389e-17 
c_198 M7:SRC M5:SRC 2.8937e-20 
c_199 M7:SRC M6:SRC 2.4313e-19 
c_200 M7:SRC M8:DRN 1.38621e-17 
c_201 M7:SRC CLK:1 5.44365e-18 
c_202 M7:SRC GND:1 3.01475e-18 
c_203 M7:SRC M8:GATE 8.84858e-18 
c_204 M7:SRC M7:GATE 1.47963e-17 
c_205 M7:SRC CLK 1.32728e-17 
c_206 M7:SRC DD1:CATHODE 5.66958e-19 
c_207 M7:SRC 0 3.83369e-18 
c_208 M3:GATE M1:SRC 4.97775e-20 
c_209 M3:GATE C 1.97379e-19 
c_210 M3:GATE M4:DRN 4.58969e-18 
c_211 M3:GATE M4:SRC 1.47697e-18 
c_212 M3:GATE GND:1 4.70252e-18 
c_213 M3:GATE M8:DRN 2.81325e-17 
c_214 M3:GATE 0 3.56505e-18 
c_215 VDD:1 CLK:1 1.13027e-17 
c_216 VDD:1 N_12:4 4.19765e-17 
c_217 VDD:1 N_12:2 2.88009e-19 
c_218 VDD:1 C 1.87559e-17 
c_219 VDD:1 M16:GATE 7.21422e-18 
c_220 VDD:1 M18:DRN 4.44775e-19 
c_221 VDD:1 M17:DRN 1.64936e-18 
c_222 VDD:1 M15:DRN 8.51175e-19 
c_223 VDD:1 M13:DRN 9.32196e-20 
c_224 VDD:1 N_12:1 2.50977e-19 
c_225 VDD:1 M11:DRN 9.32196e-20 
c_226 VDD:1 M18:GATE 1.55387e-18 
c_227 VDD:1 M15:GATE 5.74278e-18 
c_228 VDD:1 M14:GATE 1.97976e-18 
c_229 VDD:1 M13:GATE 9.23347e-19 
c_230 VDD:1 M12:GATE 3.45612e-19 
c_231 VDD:1 C:1 5.09112e-17 
c_232 VDD:1 M17:GATE 1.58933e-18 
c_233 VDD:1 0 4.13391e-17 
c_234 VDD:2 CLK:1 1.74115e-19 
c_235 VDD:2 N_12:2 1.04231e-18 
c_236 VDD:2 C 1.33458e-18 
c_237 VDD:2 M16:GATE 1.83045e-19 
c_238 VDD:2 M15:DRN 1.03413e-19 
c_239 VDD:2 M13:DRN 1.03413e-19 
c_240 VDD:2 N_12:1 9.40773e-19 
c_241 VDD:2 M11:DRN 6.30723e-20 
c_242 VDD:2 M15:GATE 3.62207e-20 
c_243 VDD:2 M14:GATE 3.03397e-19 
c_244 VDD:2 M13:GATE 4.27849e-19 
c_245 VDD:2 M12:GATE 9.80594e-19 
c_246 VDD:2 C:1 3.23531e-17 
c_247 VDD:2 M17:GATE 2.98192e-19 
c_248 VDD:2 M11:GATE 4.57012e-19 
c_249 VDD:2 M10:GATE 1.10915e-18 
c_250 VDD:2 M9:GATE 1.75137e-18 
c_251 VDD:2 0 3.52888e-17 
c_252 VDD CLK:1 3.03896e-18 
c_253 VDD N_12:4 1.56725e-16 
c_254 VDD N_12:2 7.65409e-20 
c_255 VDD C 2.02694e-17 
c_256 VDD M16:GATE 4.24801e-18 
c_257 VDD CLK 1.03479e-18 
c_258 VDD M18:DRN 1.34536e-18 
c_259 VDD M17:DRN 2.07051e-18 
c_260 VDD M15:DRN 2.64469e-18 
c_261 VDD M13:DRN 2.64469e-18 
c_262 VDD N_12:1 6.7003e-19 
c_263 VDD M11:DRN 2.64469e-18 
c_264 VDD M9:DRN 1.83749e-18 
c_265 VDD M18:GATE 3.28572e-18 
c_266 VDD M15:GATE 5.62592e-18 
c_267 VDD M14:GATE 3.28256e-18 
c_268 VDD M13:GATE 3.01967e-18 
c_269 VDD M12:GATE 3.37661e-18 
c_270 VDD C:1 9.22861e-17 
c_271 VDD M17:GATE 4.42293e-18 
c_272 VDD M11:GATE 2.84217e-18 
c_273 VDD M10:GATE 2.96076e-18 
c_274 VDD M9:GATE 6.61789e-19 
c_275 VDD 0 1.52038e-16 
c_276 M12:DRN N_12:4 7.40134e-20 
c_277 M12:DRN N_12:2 1.5982e-17 
c_278 M12:DRN C 4.96245e-18 
c_279 M12:DRN N_12:1 3.29691e-18 
c_280 M12:DRN M13:GATE 1.47201e-18 
c_281 M12:DRN M12:GATE 2.03818e-17 
c_282 M12:DRN C:1 9.41305e-18 
c_283 M12:DRN M11:GATE 1.68844e-17 
c_284 M12:DRN M10:GATE 1.52295e-18 
c_285 M12:DRN 0 6.41635e-18 
c_286 M10:DRN N_12:4 8.58205e-20 
c_287 M10:DRN N_12:2 1.48047e-17 
c_288 M10:DRN C 8.006e-18 
c_289 M10:DRN N_12:1 9.27514e-18 
c_290 M10:DRN M1:GATE 7.0857e-18 
c_291 M10:DRN C:1 2.73866e-20 
c_292 M10:DRN M11:GATE 1.45737e-18 
c_293 M10:DRN M10:GATE 2.21672e-17 
c_294 M10:DRN M9:GATE 1.41285e-17 
c_295 M10:DRN 0 4.40185e-18 
c_296 M14:DRN N_12:4 7.06552e-20 
c_297 M14:DRN N_12:2 2.85297e-18 
c_298 M14:DRN C 4.42929e-18 
c_299 M14:DRN M15:GATE 1.17145e-18 
c_300 M14:DRN M14:GATE 2.09958e-17 
c_301 M14:DRN M13:GATE 2.10065e-17 
c_302 M14:DRN M12:GATE 1.47583e-18 
c_303 M14:DRN C:1 9.233e-18 
c_304 M14:DRN 0 5.79594e-18 
c_305 M18:SRC N_12:5 1.10946e-18 
c_306 M18:SRC CLK:1 4.59252e-17 
c_307 M18:SRC N_12:4 2.81998e-17 
c_308 M18:SRC C 2.70405e-17 
c_309 M18:SRC N_12:3 1.8634e-18 
c_310 M18:SRC M16:GATE 1.32226e-17 
c_311 M18:SRC CLK 2.78176e-18 
c_312 M18:SRC M18:DRN 1.49318e-17 
c_313 M18:SRC M17:DRN 1.47202e-17 
c_314 M18:SRC M15:DRN 1.38214e-17 
c_315 M18:SRC M13:DRN 1.45146e-17 
c_316 M18:SRC N_12:1 5.76644e-18 
c_317 M18:SRC M11:DRN 1.31812e-17 
c_318 M18:SRC M9:DRN 8.62029e-18 
c_319 M18:SRC M18:GATE 4.69042e-17 
c_320 M18:SRC M15:GATE 1.10985e-17 
c_321 M18:SRC M14:GATE 1.30439e-17 
c_322 M18:SRC M13:GATE 1.41475e-17 
c_323 M18:SRC M12:GATE 1.25818e-17 
c_324 M18:SRC C:1 5.71859e-17 
c_325 M18:SRC M17:GATE 2.20857e-17 
c_326 M18:SRC M11:GATE 1.31022e-17 
c_327 M18:SRC M10:GATE 1.40464e-17 
c_328 M18:SRC M9:GATE 1.39593e-17 
c_329 M18:SRC 0 7.26569e-17 
c_330 M16:DRN CLK:1 5.25731e-18 
c_331 M16:DRN N_12:4 2.50097e-18 
c_332 M16:DRN N_12:2 4.8904e-18 
c_333 M16:DRN C 8.91649e-20 
c_334 M16:DRN M7:GATE 5.03996e-18 
c_335 M16:DRN M16:GATE 3.12393e-17 
c_336 M16:DRN M17:DRN 4.10737e-19 
c_337 M16:DRN M15:DRN 1.86833e-18 
c_338 M16:DRN M15:GATE 2.21245e-17 
c_339 M16:DRN M14:GATE 1.03096e-18 
c_340 M16:DRN C:1 2.06977e-19 
c_341 M16:DRN M17:GATE 1.1444e-18 
c_342 M16:DRN 0 9.48974e-18 

.ENDS
