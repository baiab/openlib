
.subckt INVX2  A Y
M1 GND A Y GND nch l=0.18u w=2.00u 
M2 VDD A Y VDD pch l=0.18u w=3.00u 
c_1 Y GND 8.0e-16 
c_2 A Y 2.0e-17 
c_3 A GND 8.0e-16 
.ENDS
