
.subckt ND2D1  A1 A2 ZN
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.0486p as=0.12636p l=0.09u nrd=0.167 nrs=0.433 pd=0.72u ps=1.548u sa=5.04e-07 sb=2.34e-07 w=0.54u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.12636p as=0.0486p l=0.09u nrd=0.433 nrs=0.167 pd=1.548u ps=0.72u sa=2.34e-07 sb=5.04e-07 w=0.54u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK pch ad=0.08424p as=0.16848p l=0.09u nrd=0.162 nrs=0.325 pd=0.954u ps=1.908u sa=5.58e-07 sb=2.34e-07 w=0.72u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK pch ad=0.16848p as=0.08424p l=0.09u nrd=0.325 nrs=0.162 pd=1.908u ps=0.954u sa=2.34e-07 sb=5.58e-07 w=0.72u 
R1 M1:DRN GND 18.3033
R2 M2:BULK GND 4.61359
R3 M2:BULK M1:BULK 0.001
R4 M4:DRN ZN 9.33848
R5 M4:DRN M3:SRC 0.001
R6 ZN M2:SRC 18.291
R7 M4:GATE A1 115.326
R8 M4:GATE M2:GATE 293.574
R9 A1 M2:GATE 96.7248
R10 M3:GATE A2 90.1507
R11 M3:GATE M1:GATE 275.349
R12 A2 M1:GATE 72.9533
R13 M2:DRN M1:SRC 0.001
R14 M4:BULK M3:BULK 0.001
R15 M4:BULK VDD 4.5576
R16 M4:BULK M4:SRC 1194.29
R17 VDD M3:DRN 18.2668
R18 VDD M4:SRC 18.6974
c_1 M1:DRN 0 3.62051e-18 
c_2 M2:BULK 0 2.74534e-17 
c_3 GND 0 7.72146e-17 
c_4 M4:DRN GND 3.87767e-19 
c_5 M4:DRN M2:BULK 6.72634e-19 
c_6 M4:DRN 0 5.60204e-18 
c_7 ZN GND 4.22304e-17 
c_8 ZN M1:DRN 7.55283e-20 
c_9 ZN M2:BULK 9.47618e-18 
c_10 ZN 0 1.76191e-17 
c_11 M2:SRC M2:BULK 8.97676e-18 
c_12 M2:SRC M1:DRN 1.45997e-18 
c_13 M2:SRC GND 1.74936e-18 
c_14 M2:SRC 0 2.61256e-18 
c_15 M4:GATE M4:DRN 3.34301e-17 
c_16 M4:GATE ZN 1.0976e-17 
c_17 M4:GATE 0 7.65839e-18 
c_18 A1 GND 7.26207e-18 
c_19 A1 M1:DRN 2.48449e-19 
c_20 A1 M4:DRN 2.92691e-18 
c_21 A1 ZN 1.14973e-16 
c_22 A1 M2:BULK 1.15078e-17 
c_23 A1 M2:SRC 6.33396e-19 
c_24 A1 0 1.019e-17 
c_25 M2:GATE M2:BULK 1.60755e-17 
c_26 M2:GATE ZN 1.59611e-18 
c_27 M2:GATE M2:SRC 3.19572e-17 
c_28 M2:GATE GND 9.25502e-18 
c_29 M2:GATE 0 9.10836e-18 
c_30 M3:GATE M4:GATE 1.16163e-17 
c_31 M3:GATE M4:DRN 3.5177e-17 
c_32 M3:GATE ZN 8.51038e-18 
c_33 M3:GATE M2:BULK 2.12664e-18 
c_34 M3:GATE 0 1.63354e-17 
c_35 A2 GND 3.69234e-17 
c_36 A2 M1:DRN 3.23021e-17 
c_37 A2 M4:DRN 1.86847e-18 
c_38 A2 ZN 3.5829e-17 
c_39 A2 M2:BULK 4.54625e-18 
c_40 A2 A1 2.03602e-17 
c_41 A2 M4:GATE 2.37908e-19 
c_42 A2 0 5.3127e-19 
c_43 M1:GATE ZN 8.28407e-18 
c_44 M1:GATE A1 1.10109e-17 
c_45 M1:GATE M2:BULK 2.14002e-17 
c_46 M1:GATE M2:GATE 6.95408e-18 
c_47 M1:GATE M2:SRC 1.60689e-19 
c_48 M1:GATE GND 6.59538e-18 
c_49 M1:GATE 0 1.02796e-17 
c_50 M2:DRN M4:DRN 3.52868e-18 
c_51 M2:DRN ZN 7.30478e-19 
c_52 M2:DRN M2:BULK 6.53071e-18 
c_53 M2:DRN GND 5.10278e-19 
c_54 M2:DRN 0 1.21796e-19 
c_55 M4:BULK M3:GATE 1.67917e-17 
c_56 M4:BULK M4:GATE 1.67902e-17 
c_57 M4:BULK M4:DRN 1.34705e-17 
c_58 M4:BULK ZN 8.14285e-18 
c_59 M4:BULK A2 1.00353e-17 
c_60 M4:BULK A1 1.1488e-17 
c_61 M4:BULK 0 2.88464e-17 
c_62 VDD M3:GATE 1.55179e-17 
c_63 VDD M4:GATE 1.49379e-17 
c_64 VDD M4:DRN 3.04627e-18 
c_65 VDD ZN 9.64169e-17 
c_66 VDD A2 2.10702e-17 
c_67 VDD A1 1.50479e-17 
c_68 VDD 0 8.62357e-17 
c_69 M3:DRN M4:GATE 2.09883e-20 
c_70 M3:DRN M3:GATE 1.66998e-17 
c_71 M3:DRN M4:DRN 2.77945e-19 
c_72 M3:DRN ZN 5.79208e-19 
c_73 M3:DRN A2 1.63131e-17 
c_74 M3:DRN 0 2.68442e-18 
c_75 M4:SRC M4:DRN 2.77945e-19 
c_76 M4:SRC M4:GATE 3.03118e-17 
c_77 M4:SRC M3:GATE 2.09883e-20 
c_78 M4:SRC ZN 1.00756e-18 
c_79 M4:SRC A1 2.74379e-18 
c_80 M4:SRC M2:SRC 2.08295e-18 
c_81 M4:SRC 0 8.42058e-19 

.ENDS
