
.subckt AOI33D4  A1 A2 A3 B1 B2 B3 ZN
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=2.412e-06 sb=1.116e-06 w=0.54u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.06318p as=0.07371p l=0.09u nrd=0.217 nrs=0.254 pd=0.774u ps=0.963u sa=2.088e-06 sb=1.44e-06 w=0.54u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.05103p as=0.05103p l=0.09u nrd=0.175 nrs=0.175 pd=0.729u ps=0.729u sa=1.494e-06 sb=2.034e-06 w=0.54u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.0486p as=0.0486p l=0.09u nrd=0.167 nrs=0.167 pd=0.72u ps=0.72u sa=5.04e-07 sb=3.024e-06 w=0.54u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.05103p as=0.09477p l=0.09u nrd=0.175 nrs=0.325 pd=0.729u ps=0.891u sa=1.215e-06 sb=2.313e-06 w=0.54u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=2.691e-06 sb=8.37e-07 w=0.54u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.06075p as=0.12636p l=0.09u nrd=0.209 nrs=0.433 pd=0.927u ps=1.548u sa=3.294e-06 sb=2.34e-07 w=0.54u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.05103p as=0.07371p l=0.09u nrd=0.175 nrs=0.254 pd=0.729u ps=0.963u sa=1.773e-06 sb=1.755e-06 w=0.54u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.12636p as=0.0486p l=0.09u nrd=0.433 nrs=0.167 pd=1.548u ps=0.72u sa=2.34e-07 sb=3.294e-06 w=0.54u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.0486p as=0.09477p l=0.09u nrd=0.167 nrs=0.325 pd=0.72u ps=0.891u sa=7.74e-07 sb=2.754e-06 w=0.54u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=3.015e-06 sb=5.13e-07 w=0.54u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK pch ad=0.08424p as=0.08181p l=0.09u nrd=0.162 nrs=0.158 pd=0.954u ps=1.116u sa=1.836e-06 sb=1.728e-06 w=0.72u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=2.727e-06 sb=8.37e-07 w=0.72u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK pch ad=0.16848p as=0.09072p l=0.09u nrd=0.325 nrs=0.175 pd=1.908u ps=0.972u sa=2.34e-07 sb=3.33e-06 w=0.72u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK pch ad=0.08424p as=0.08424p l=0.09u nrd=0.162 nrs=0.162 pd=0.954u ps=0.954u sa=9e-07 sb=2.664e-06 w=0.72u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=2.448e-06 sb=1.116e-06 w=0.72u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=3.051e-06 sb=5.13e-07 w=0.72u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK pch ad=0.08424p as=0.08181p l=0.09u nrd=0.162 nrs=0.158 pd=0.954u ps=1.116u sa=1.512e-06 sb=2.052e-06 w=0.72u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK pch ad=0.07776p as=0.16848p l=0.09u nrd=0.15 nrs=0.325 pd=1.107u ps=1.908u sa=3.33e-06 sb=2.34e-07 w=0.72u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK pch ad=0.09072p as=0.08424p l=0.09u nrd=0.175 nrs=0.162 pd=0.972u ps=0.954u sa=5.76e-07 sb=2.988e-06 w=0.72u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK pch ad=0.08424p as=0.08181p l=0.09u nrd=0.162 nrs=0.158 pd=0.954u ps=1.116u sa=1.224e-06 sb=2.34e-06 w=0.72u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK pch ad=0.08424p as=0.08181p l=0.09u nrd=0.162 nrs=0.158 pd=0.954u ps=1.116u sa=2.124e-06 sb=1.44e-06 w=0.72u 
R1 M1:DRN M2:DRN 0.001
R2 M2:SRC M6:DRN 0.001
R3 M5:DRN M4:SRC 0.001
R4 M4:DRN M3:SRC 0.001
R5 M15:DRN M17:DRN 54.487
R6 M15:DRN M12:DRN 55.7852
R7 M15:DRN M14:SRC 0.001
R8 M17:DRN M12:DRN 54.4002
R9 M17:DRN M16:SRC 0.001
R10 M12:DRN M13:DRN 0.001
R11 M12:GATE B3 97.6288
R12 M12:GATE M1:GATE 310.85
R13 B3 M1:GATE 74.1531
R14 M13:GATE B2 93.9105
R15 M13:GATE M2:GATE 313.473
R16 B2 M2:GATE 77.4391
R17 M17:GATE M6:GATE 297.009
R18 M17:GATE B1 92.3837
R19 B1 M6:GATE 75.4797
R20 M16:GATE A1 97.0066
R21 M16:GATE M5:GATE 303.137
R22 A1 M5:GATE 73.3876
R23 M15:GATE M4:GATE 305.443
R24 M15:GATE A2 93.2367
R25 A2 M4:GATE 76.4373
R26 M14:GATE A3 115.326
R27 M14:GATE M3:GATE 293.574
R28 A3 M3:GATE 96.7248
R29 M10:BULK M1:SRC 1.4735e-05
R30 M10:BULK M3:BULK 0.001
R31 M10:BULK M4:BULK 0.001
R32 M10:BULK M5:BULK 0.001
R33 M10:BULK M6:BULK 0.001
R34 M10:BULK M2:BULK 0.001
R35 M10:BULK M1:BULK 0.001
R36 M10:BULK M9:BULK 0.001
R37 M10:BULK M8:BULK 0.001
R38 M10:BULK M7:BULK 0.001
R39 M10:BULK M11:BULK 0.001
R40 M9:DRN M8:SRC 0.001
R41 M9:DRN M1:SRC 2e-09
R42 M7:SRC M11:DRN 0.001
R43 M7:SRC M1:SRC 2e-09
R44 GND M1:SRC 1.38966
R45 GND M3:DRN 18.1744
R46 M1:SRC M10:SRC 0.001
R47 ZN M10:DRN 18.2086
R48 ZN M19:DRN 9.3497
R49 ZN M21:DRN 9.37828
R50 ZN M7:DRN 18.1975
R51 M21:DRN M20:DRN 0.001
R52 M21:DRN M19:DRN 608.583
R53 M7:DRN M8:DRN 0.001
R54 M19:DRN M18:DRN 0.001
R55 M10:DRN M9:SRC 0.001
R56 M19:BULK M21:BULK 0.001
R57 M19:BULK M17:SRC 1.46592e-05
R58 M19:BULK M12:SRC 0.00514403
R59 M19:BULK M18:SRC 0.00561167
R60 M19:BULK M20:SRC 0.00561167
R61 M19:BULK M20:BULK 0.001
R62 M19:BULK M22:BULK 0.001
R63 M19:BULK M14:BULK 0.001
R64 M19:BULK M15:BULK 0.001
R65 M19:BULK M16:BULK 0.001
R66 M19:BULK M17:BULK 0.001
R67 M19:BULK M13:BULK 0.001
R68 M19:BULK M12:BULK 0.001
R69 M19:BULK M18:BULK 0.001
R70 VDD M17:SRC 2.83169
R71 VDD M18:SRC 50.2227
R72 VDD VDD:1 0.602257
R73 VDD:1 M18:SRC 7.01922
R74 VDD:1 M20:SRC 9.01083
R75 VDD:1 M17:SRC 5.46238
R76 M18:SRC M17:SRC 1.52222e-09
R77 M18:SRC M20:SRC 1.12222e-09
R78 M18:SRC M21:SRC 0.001
R79 M20:SRC M22:DRN 0.001
R80 M17:SRC M12:SRC 7.22222e-10
R81 M17:SRC M13:SRC 0.001
R82 M12:SRC M19:SRC 0.001
R83 N_4:1 N_4:2 35.4222
R84 N_4:1 M20:GATE 66.96
R85 N_4:1 M8:GATE 130.719
R86 N_4:1 M7:GATE 47.5765
R87 N_4:1 M11:SRC 66.4936
R88 N_4:1 M22:SRC 32.3266
R89 N_4:1 M21:GATE 155.858
R90 N_4:2 M10:GATE 88.655
R91 N_4:2 M19:GATE 105.704
R92 N_4:2 M9:GATE 44.28
R93 N_4:2 M8:GATE 147.519
R94 N_4:2 M18:GATE 55.08
R95 N_4:2 M21:GATE 175.889
R96 M22:SRC M11:SRC 38.3222
R97 M21:GATE M8:GATE 649.086
R98 M19:GATE M10:GATE 335.904
R99 N_9:1 M6:SRC 64.4112
R100 N_9:1 M14:DRN 74.2796
R101 N_9:1 M16:DRN 75.1363
R102 N_9:1 M11:GATE 47.1388
R103 N_9:1 M22:GATE 64.4188
R104 M16:DRN M6:SRC 79.3911
R105 M16:DRN M14:DRN 69.6472
R106 M16:DRN M15:SRC 0.001
R107 M14:DRN M6:SRC 78.4858
R108 M6:SRC M5:SRC 0.001
c_1 M1:DRN 0 1.93948e-19 
c_2 M2:SRC 0 9.03394e-20 
c_3 M5:DRN 0 4.34055e-20 
c_4 M4:DRN 0 1.20977e-19 
c_5 M15:DRN M4:DRN 3.4991e-18 
c_6 M15:DRN 0 2.11943e-17 
c_7 M17:DRN 0 2.48075e-19 
c_8 M12:DRN M1:DRN 3.81856e-18 
c_9 M12:DRN 0 3.69715e-18 
c_10 M12:GATE M15:DRN 5.92997e-18 
c_11 M12:GATE M12:DRN 1.68709e-17 
c_12 M12:GATE 0 5.36327e-18 
c_13 B3 M15:DRN 1.09028e-17 
c_14 B3 M12:DRN 4.43971e-18 
c_15 B3 0 5.10184e-18 
c_16 M1:GATE 0 2.54576e-18 
c_17 M13:GATE M12:GATE 1.12683e-17 
c_18 M13:GATE B3 4.38109e-18 
c_19 M13:GATE M17:DRN 1.36697e-19 
c_20 M13:GATE M12:DRN 2.91473e-17 
c_21 M13:GATE 0 7.96852e-18 
c_22 B2 M12:GATE 1.51774e-18 
c_23 B2 M1:DRN 2.89307e-18 
c_24 B2 B3 9.09705e-17 
c_25 B2 M2:SRC 1.94388e-18 
c_26 B2 M12:DRN 1.23654e-17 
c_27 B2 0 4.91459e-18 
c_28 M2:GATE M12:DRN 1.24134e-19 
c_29 M2:GATE B3 2.59077e-17 
c_30 M2:GATE M1:GATE 6.09739e-18 
c_31 M2:GATE 0 3.93875e-18 
c_32 M17:GATE M17:DRN 1.6586e-17 
c_33 M17:GATE B2 8.18661e-18 
c_34 M17:GATE M12:DRN 8.01345e-18 
c_35 M17:GATE M13:GATE 1.71549e-17 
c_36 M17:GATE 0 9.62795e-18 
c_37 B1 M2:SRC 3.02517e-18 
c_38 B1 M17:DRN 3.13271e-18 
c_39 B1 B2 7.7616e-17 
c_40 B1 M12:DRN 1.52025e-17 
c_41 B1 M13:GATE 2.15386e-18 
c_42 B1 0 9.17702e-18 
c_43 M6:GATE B2 2.71604e-17 
c_44 M6:GATE M2:GATE 6.44501e-18 
c_45 M6:GATE 0 1.19992e-18 
c_46 M16:GATE M15:DRN 1.06341e-19 
c_47 M16:GATE M17:DRN 1.67375e-17 
c_48 M16:GATE M17:GATE 1.1832e-17 
c_49 M16:GATE B1 1.94678e-18 
c_50 M16:GATE M12:DRN 6.72632e-18 
c_51 M16:GATE 0 5.60844e-18 
c_52 A1 M17:DRN 7.10361e-19 
c_53 A1 M17:GATE 5.14677e-20 
c_54 A1 B1 6.10852e-17 
c_55 A1 M12:DRN 5.05162e-18 
c_56 A1 0 2.89152e-18 
c_57 M5:GATE B1 1.79877e-17 
c_58 M5:GATE M6:GATE 3.3212e-18 
c_59 M5:GATE 0 1.08261e-18 
c_60 M15:GATE M15:DRN 1.66051e-17 
c_61 M15:GATE A1 7.44497e-18 
c_62 M15:GATE M16:GATE 1.19152e-17 
c_63 M15:GATE M17:DRN 1.06341e-19 
c_64 M15:GATE M12:DRN 6.83276e-18 
c_65 M15:GATE 0 7.6999e-18 
c_66 A2 M4:DRN 2.83756e-18 
c_67 A2 M15:DRN 8.15015e-18 
c_68 A2 M5:DRN 2.98041e-18 
c_69 A2 A1 5.18879e-17 
c_70 A2 M16:GATE 1.44264e-18 
c_71 A2 M12:DRN 1.41449e-18 
c_72 A2 0 5.53947e-18 
c_73 M4:GATE A1 2.80054e-17 
c_74 M4:GATE M5:GATE 7.15092e-18 
c_75 M4:GATE 0 6.14076e-19 
c_76 M14:GATE M15:DRN 1.31793e-17 
c_77 M14:GATE M15:GATE 1.00431e-17 
c_78 M14:GATE M12:DRN 4.43865e-18 
c_79 M14:GATE A2 1.40663e-18 
c_80 M14:GATE 0 2.33464e-17 
c_81 A3 M15:DRN 2.77243e-18 
c_82 A3 M15:GATE 9.83486e-20 
c_83 A3 M17:DRN 2.29681e-19 
c_84 A3 A2 3.87596e-17 
c_85 A3 0 1.33373e-18 
c_86 M3:GATE A2 2.49647e-19 
c_87 M3:GATE M4:GATE 6.84796e-18 
c_88 M3:GATE 0 3.94867e-18 
c_89 M10:BULK M12:GATE 2.88614e-18 
c_90 M10:BULK B3 2.60902e-18 
c_91 M10:BULK M1:GATE 3.94486e-18 
c_92 M10:BULK A3 4.87366e-18 
c_93 M10:BULK M3:GATE 9.05714e-18 
c_94 M10:BULK M4:GATE 4.74693e-18 
c_95 M10:BULK M15:GATE 2.60632e-18 
c_96 M10:BULK A1 2.90556e-18 
c_97 M10:BULK M5:GATE 4.8575e-18 
c_98 M10:BULK M16:GATE 4.21817e-18 
c_99 M10:BULK M17:GATE 2.2574e-18 
c_100 M10:BULK M6:GATE 5.65277e-18 
c_101 M10:BULK B1 9.05904e-19 
c_102 M10:BULK B2 2.94261e-18 
c_103 M10:BULK M2:GATE 3.5057e-18 
c_104 M10:BULK A2 1.12252e-18 
c_105 M10:BULK M13:GATE 2.95346e-18 
c_106 M9:DRN 0 2.7552e-18 
c_107 M7:SRC 0 2.97259e-18 
c_108 GND M1:DRN 3.71476e-19 
c_109 GND B3 2.38653e-18 
c_110 GND M1:GATE 4.75254e-18 
c_111 GND M2:SRC 3.71476e-19 
c_112 GND A3 1.50509e-17 
c_113 GND M3:GATE 6.61983e-18 
c_114 GND M4:DRN 4.77015e-19 
c_115 GND M4:GATE 6.57206e-18 
c_116 GND M5:DRN 3.71476e-19 
c_117 GND A1 3.06723e-18 
c_118 GND M5:GATE 7.20443e-18 
c_119 GND M6:GATE 4.93921e-18 
c_120 GND B1 2.05258e-18 
c_121 GND B2 1.91439e-18 
c_122 GND M2:GATE 4.82231e-18 
c_123 GND A2 1.3841e-18 
c_124 GND 0 1.43019e-16 
c_125 M3:DRN A2 1.71014e-19 
c_126 M3:DRN M3:GATE 1.67807e-17 
c_127 M3:DRN A3 1.81401e-17 
c_128 M3:DRN M5:DRN 7.51687e-19 
c_129 M1:SRC M1:DRN 6.84748e-18 
c_130 M1:SRC B3 1.79534e-18 
c_131 M1:SRC M1:GATE 2.52284e-17 
c_132 M1:SRC M2:SRC 6.92586e-18 
c_133 M1:SRC A3 6.65229e-19 
c_134 M1:SRC M3:GATE 9.4396e-18 
c_135 M1:SRC M4:DRN 6.52898e-18 
c_136 M1:SRC M4:GATE 9.44127e-18 
c_137 M1:SRC M15:GATE 2.68077e-19 
c_138 M1:SRC M5:DRN 6.53001e-18 
c_139 M1:SRC A1 4.509e-19 
c_140 M1:SRC M5:GATE 9.44066e-18 
c_141 M1:SRC M16:GATE 2.83352e-19 
c_142 M1:SRC M17:GATE 4.06848e-19 
c_143 M1:SRC M6:GATE 9.44138e-18 
c_144 M1:SRC B1 5.59607e-19 
c_145 M1:SRC B2 6.18578e-19 
c_146 M1:SRC M2:GATE 1.13508e-17 
c_147 M1:SRC 0 1.10264e-16 
c_148 ZN M1:SRC 2.27494e-18 
c_149 ZN M12:GATE 3.67071e-18 
c_150 ZN GND 5.15011e-18 
c_151 ZN B3 2.74368e-17 
c_152 ZN M1:GATE 8.82884e-19 
c_153 ZN M10:BULK 5.58554e-19 
c_154 ZN M9:DRN 3.35989e-18 
c_155 ZN 0 1.87199e-17 
c_156 M21:DRN M1:SRC 4.42193e-20 
c_157 M21:DRN 0 3.46972e-18 
c_158 M7:DRN M1:SRC 8.82966e-18 
c_159 M7:DRN GND 1.34188e-18 
c_160 M7:DRN 0 1.49171e-18 
c_161 M19:DRN M1:SRC 1.81772e-20 
c_162 M19:DRN M12:GATE 4.89297e-19 
c_163 M19:DRN 0 3.63686e-18 
c_164 M10:DRN M1:SRC 8.44104e-18 
c_165 M10:DRN GND 1.30149e-18 
c_166 M10:DRN B3 1.00655e-19 
c_167 M10:DRN M1:GATE 3.60467e-19 
c_168 M10:DRN 0 1.52113e-18 
c_169 M19:BULK M12:GATE 7.36708e-18 
c_170 M19:BULK B3 3.63438e-18 
c_171 M19:BULK ZN 1.23795e-17 
c_172 M19:BULK A3 6.50447e-18 
c_173 M19:BULK M15:DRN 9.21939e-18 
c_174 M19:BULK M15:GATE 8.61537e-18 
c_175 M19:BULK M5:DRN 4.60357e-19 
c_176 M19:BULK A1 2.71805e-18 
c_177 M19:BULK M16:GATE 7.3468e-18 
c_178 M19:BULK M17:GATE 6.55066e-18 
c_179 M19:BULK B1 2.77762e-18 
c_180 M19:BULK B2 4.77268e-18 
c_181 M19:BULK M19:DRN 5.14489e-18 
c_182 M19:BULK M21:DRN 1.7583e-18 
c_183 M19:BULK A2 9.99315e-19 
c_184 M19:BULK M13:GATE 7.17228e-18 
c_185 M19:BULK M14:GATE 6.87973e-18 
c_186 VDD M12:GATE 7.48509e-18 
c_187 VDD B3 3.10741e-18 
c_188 VDD ZN 9.46939e-17 
c_189 VDD A3 1.08917e-18 
c_190 VDD M15:DRN 2.93197e-18 
c_191 VDD M15:GATE 8.27999e-18 
c_192 VDD M16:GATE 8.2635e-18 
c_193 VDD M17:DRN 1.34489e-16 
c_194 VDD M17:GATE 7.57721e-18 
c_195 VDD B1 7.74334e-19 
c_196 VDD B2 9.1311e-20 
c_197 VDD M12:DRN 4.9906e-17 
c_198 VDD M19:DRN 2.67113e-18 
c_199 VDD M21:DRN 2.76019e-18 
c_200 VDD M13:GATE 7.44826e-18 
c_201 VDD M14:GATE 9.51135e-18 
c_202 VDD 0 1.30476e-16 
c_203 VDD:1 0 7.90364e-18 
c_204 M18:SRC ZN 1.36331e-17 
c_205 M18:SRC M21:DRN 1.07984e-18 
c_206 M18:SRC 0 5.91481e-18 
c_207 M20:SRC ZN 1.04817e-19 
c_208 M20:SRC 0 6.71293e-18 
c_209 M17:SRC M10:DRN 8.11934e-21 
c_210 M17:SRC M12:GATE 1.03312e-17 
c_211 M17:SRC B3 5.84627e-19 
c_212 M17:SRC ZN 7.02861e-19 
c_213 M17:SRC M2:SRC 3.09066e-18 
c_214 M17:SRC A3 3.62231e-19 
c_215 M17:SRC M15:DRN 1.2111e-17 
c_216 M17:SRC M15:GATE 9.51257e-18 
c_217 M17:SRC M5:DRN 2.67452e-19 
c_218 M17:SRC A1 2.05808e-20 
c_219 M17:SRC M16:GATE 1.01848e-17 
c_220 M17:SRC M17:DRN 1.14747e-17 
c_221 M17:SRC M17:GATE 1.97445e-17 
c_222 M17:SRC B1 7.69871e-18 
c_223 M17:SRC B2 1.01989e-18 
c_224 M17:SRC M12:DRN 1.9235e-17 
c_225 M17:SRC M19:DRN 1.11007e-17 
c_226 M17:SRC M21:DRN 1.02793e-17 
c_227 M17:SRC M7:DRN 3.81007e-20 
c_228 M17:SRC M13:GATE 1.9816e-17 
c_229 M17:SRC M14:GATE 9.49826e-18 
c_230 M17:SRC 0 9.95051e-17 
c_231 M12:SRC M12:GATE 1.03177e-17 
c_232 M12:SRC B3 3.87862e-18 
c_233 M12:SRC ZN 4.87043e-19 
c_234 M12:SRC M12:DRN 2.74163e-21 
c_235 M12:SRC M13:GATE 8.3293e-19 
c_236 M12:SRC 0 3.53833e-18 
c_237 N_4:1 M10:DRN 1.47635e-19 
c_238 N_4:1 M1:SRC 1.31919e-19 
c_239 N_4:1 GND 1.33082e-18 
c_240 N_4:1 M17:SRC 6.5796e-21 
c_241 N_4:1 M10:BULK 8.44771e-19 
c_242 N_4:1 M19:BULK 6.92212e-18 
c_243 N_4:1 ZN 1.20237e-16 
c_244 N_4:1 VDD 7.76493e-21 
c_245 N_4:1 M18:SRC 8.4926e-21 
c_246 N_4:1 M21:DRN 2.83788e-18 
c_247 N_4:1 M7:DRN 2.41016e-17 
c_248 N_4:1 M7:SRC 2.18325e-19 
c_249 N_4:1 0 1.07893e-21 
c_250 N_4:2 M10:DRN 3.00057e-17 
c_251 N_4:2 M1:SRC 5.45316e-19 
c_252 N_4:2 M12:GATE 3.31223e-18 
c_253 N_4:2 GND 1.26081e-18 
c_254 N_4:2 M17:SRC 7.88775e-20 
c_255 N_4:2 B3 9.30965e-18 
c_256 N_4:2 M1:GATE 1.65308e-17 
c_257 N_4:2 M10:BULK 7.67655e-18 
c_258 N_4:2 M19:BULK 3.56992e-18 
c_259 N_4:2 ZN 3.67515e-17 
c_260 N_4:2 VDD 5.70019e-19 
c_261 N_4:2 M19:DRN 1.42589e-17 
c_262 N_4:2 M9:DRN 9.38217e-18 
c_263 N_4:2 M18:SRC 9.78363e-18 
c_264 N_4:2 M21:DRN 1.404e-17 
c_265 N_4:2 M7:DRN 9.65567e-18 
c_266 N_4:2 0 9.70945e-19 
c_267 M22:SRC M1:SRC 8.85342e-19 
c_268 M22:SRC M12:GATE 1.81621e-19 
c_269 M22:SRC GND 1.8735e-17 
c_270 M22:SRC M17:SRC 9.99791e-18 
c_271 M22:SRC B3 1.23163e-18 
c_272 M22:SRC M10:BULK 4.96145e-18 
c_273 M22:SRC M19:BULK 3.73081e-18 
c_274 M22:SRC VDD 3.99089e-17 
c_275 M22:SRC M19:DRN 1.39646e-20 
c_276 M22:SRC M18:SRC 2.35214e-19 
c_277 M22:SRC M21:DRN 6.57189e-19 
c_278 M22:SRC M20:SRC 5.81719e-19 
c_279 M22:SRC 0 1.36691e-18 
c_280 M21:GATE M17:SRC 4.35799e-18 
c_281 M21:GATE M19:BULK 4.3025e-18 
c_282 M21:GATE ZN 1.76717e-17 
c_283 M21:GATE VDD 7.87727e-18 
c_284 M21:GATE M19:DRN 2.95269e-19 
c_285 M21:GATE M18:SRC 1.52327e-17 
c_286 M21:GATE M21:DRN 3.52213e-17 
c_287 M21:GATE M7:DRN 2.44473e-18 
c_288 M21:GATE M20:SRC 8.3293e-19 
c_289 M21:GATE 0 2.70542e-18 
c_290 M20:GATE M20:SRC 1.00916e-17 
c_291 M20:GATE ZN 6.25388e-18 
c_292 M20:GATE M18:SRC 5.97408e-18 
c_293 M20:GATE M19:BULK 6.29979e-18 
c_294 M20:GATE VDD 7.8635e-18 
c_295 M20:GATE M21:DRN 3.3852e-17 
c_296 M20:GATE M17:SRC 4.35799e-18 
c_297 M20:GATE 0 7.97026e-19 
c_298 M7:GATE ZN 1.12647e-19 
c_299 M7:GATE M10:BULK 4.66096e-18 
c_300 M7:GATE M9:DRN 1.53101e-18 
c_301 M7:GATE M7:SRC 1.00916e-17 
c_302 M7:GATE GND 4.62058e-18 
c_303 M7:GATE M1:SRC 9.44169e-18 
c_304 M8:GATE M1:SRC 9.44169e-18 
c_305 M8:GATE GND 5.08966e-18 
c_306 M8:GATE M10:BULK 4.68688e-18 
c_307 M8:GATE ZN 1.40809e-19 
c_308 M8:GATE M9:DRN 1.00263e-17 
c_309 M8:GATE M7:DRN 1.32899e-17 
c_310 M8:GATE M7:SRC 8.3293e-19 
c_311 M11:SRC M1:SRC 9.35222e-18 
c_312 M11:SRC GND 1.78012e-18 
c_313 M11:SRC M17:SRC 3.06117e-20 
c_314 M11:SRC M7:DRN 7.51687e-19 
c_315 M11:SRC M20:SRC 4.49768e-18 
c_316 M11:SRC 0 5.35887e-17 
c_317 M19:GATE M10:DRN 5.78553e-18 
c_318 M19:GATE M12:GATE 1.79473e-17 
c_319 M19:GATE M17:SRC 9.11612e-18 
c_320 M19:GATE B3 1.8693e-18 
c_321 M19:GATE M19:BULK 4.96134e-18 
c_322 M19:GATE ZN 1.22873e-17 
c_323 M19:GATE VDD 7.89851e-18 
c_324 M19:GATE M12:SRC 1.03177e-17 
c_325 M19:GATE M19:DRN 3.37041e-17 
c_326 M19:GATE M18:SRC 8.3293e-19 
c_327 M19:GATE 0 1.96918e-18 
c_328 M18:GATE M12:GATE 1.42323e-19 
c_329 M18:GATE M17:SRC 5.17457e-18 
c_330 M18:GATE B3 2.05233e-19 
c_331 M18:GATE M19:BULK 3.68952e-18 
c_332 M18:GATE ZN 2.03525e-17 
c_333 M18:GATE VDD 8.09945e-18 
c_334 M18:GATE M12:SRC 8.3293e-19 
c_335 M18:GATE M19:DRN 3.33164e-17 
c_336 M18:GATE M18:SRC 1.40331e-17 
c_337 M18:GATE M21:DRN 2.95269e-19 
c_338 M18:GATE 0 2.0932e-18 
c_339 M10:GATE M10:DRN 1.28345e-17 
c_340 M10:GATE M1:SRC 2.00865e-17 
c_341 M10:GATE M12:GATE 3.9153e-18 
c_342 M10:GATE GND 5.35911e-18 
c_343 M10:GATE M1:GATE 3.40576e-18 
c_344 M10:GATE M10:BULK 5.08477e-18 
c_345 M10:GATE M19:BULK 3.24448e-19 
c_346 M10:GATE ZN 6.34468e-18 
c_347 M10:GATE M9:DRN 8.3293e-19 
c_348 M10:GATE 0 3.89545e-19 
c_349 M9:GATE M7:DRN 1.47635e-19 
c_350 M9:GATE ZN 6.30647e-18 
c_351 M9:GATE M9:DRN 1.00916e-17 
c_352 M9:GATE M10:BULK 4.07579e-18 
c_353 M9:GATE GND 4.87188e-18 
c_354 M9:GATE M1:GATE 2.51872e-19 
c_355 M9:GATE M1:SRC 1.06032e-17 
c_356 M9:GATE M10:DRN 9.71705e-19 
c_357 M9:GATE 0 7.5362e-19 
c_358 N_9:1 M1:SRC 1.87767e-19 
c_359 N_9:1 M12:GATE 1.24231e-20 
c_360 N_9:1 GND 3.11828e-16 
c_361 N_9:1 M17:SRC 5.48497e-20 
c_362 N_9:1 B3 9.64427e-22 
c_363 N_9:1 N_4:2 1.19365e-17 
c_364 N_9:1 M10:BULK 5.6848e-18 
c_365 N_9:1 M19:BULK 4.02241e-18 
c_366 N_9:1 ZN 2.53583e-19 
c_367 N_9:1 N_4:1 8.29419e-18 
c_368 N_9:1 VDD 6.10191e-19 
c_369 N_9:1 M5:GATE 3.49057e-19 
c_370 N_9:1 M17:DRN 4.67195e-19 
c_371 N_9:1 M8:GATE 3.0614e-19 
c_372 N_9:1 M7:DRN 1.47635e-19 
c_373 N_9:1 M7:GATE 1.01052e-17 
c_374 N_9:1 M7:SRC 3.72969e-18 
c_375 N_9:1 M20:SRC 1.43197e-19 
c_376 N_9:1 M11:SRC 3.2118e-17 
c_377 N_9:1 M22:SRC 1.92598e-20 
c_378 N_9:1 M3:DRN 1.34393e-18 
c_379 N_9:1 M13:GATE 4.19523e-19 
c_380 N_9:1 M14:GATE 1.13315e-17 
c_381 N_9:1 M21:GATE 2.0332e-18 
c_382 N_9:1 0 4.02484e-20 
c_383 M22:GATE M17:SRC 4.35799e-18 
c_384 M22:GATE M19:BULK 3.05999e-18 
c_385 M22:GATE ZN 2.47449e-18 
c_386 M22:GATE M20:GATE 1.89097e-17 
c_387 M22:GATE VDD 9.58684e-18 
c_388 M22:GATE M15:DRN 5.13037e-19 
c_389 M22:GATE M21:DRN 2.95269e-19 
c_390 M22:GATE M20:SRC 1.88127e-17 
c_391 M22:GATE M11:SRC 1.11731e-17 
c_392 M22:GATE M22:SRC 3.39994e-17 
c_393 M22:GATE M21:GATE 1.52009e-19 
c_394 M22:GATE 0 6.66343e-18 
c_395 M16:DRN M1:SRC 5.56631e-19 
c_396 M16:DRN M17:SRC 8.99778e-18 
c_397 M16:DRN M10:BULK 2.16417e-17 
c_398 M16:DRN ZN 1.18715e-16 
c_399 M16:DRN N_4:1 4.63783e-18 
c_400 M16:DRN VDD 1.27808e-18 
c_401 M16:DRN M15:GATE 1.73855e-17 
c_402 M16:DRN M5:DRN 3.00881e-18 
c_403 M16:DRN A1 8.08022e-18 
c_404 M16:DRN M16:GATE 1.67445e-17 
c_405 M16:DRN M17:GATE 3.12375e-19 
c_406 M16:DRN B1 6.68176e-20 
c_407 M16:DRN M12:DRN 5.88022e-18 
c_408 M16:DRN M7:DRN 5.96326e-18 
c_409 M16:DRN M7:SRC 3.73098e-18 
c_410 M16:DRN M22:SRC 1.26136e-16 
c_411 M16:DRN A2 9.7241e-19 
c_412 M16:DRN M14:GATE 9.00782e-20 
c_413 M16:DRN 0 1.24552e-17 
c_414 M11:GATE M7:GATE 3.85167e-18 
c_415 M11:GATE M8:GATE 2.12819e-19 
c_416 M11:GATE M10:BULK 3.81748e-18 
c_417 M11:GATE M7:SRC 1.08666e-17 
c_418 M11:GATE M11:SRC 1.23711e-17 
c_419 M11:GATE GND 6.4322e-18 
c_420 M11:GATE M1:SRC 9.44169e-18 
c_421 M11:GATE 0 1.72574e-18 
c_422 M14:DRN M1:SRC 1.47353e-17 
c_423 M14:DRN M17:SRC 9.01211e-18 
c_424 M14:DRN B3 2.6271e-17 
c_425 M14:DRN N_4:2 1.11742e-17 
c_426 M14:DRN M19:BULK 1.03215e-17 
c_427 M14:DRN M9:GATE 4.3572e-19 
c_428 M14:DRN ZN 1.33376e-17 
c_429 M14:DRN N_4:1 1.41924e-17 
c_430 M14:DRN A3 1.90446e-17 
c_431 M14:DRN VDD 1.30502e-18 
c_432 M14:DRN M15:DRN 9.70074e-17 
c_433 M14:DRN M15:GATE 9.00782e-20 
c_434 M14:DRN A1 5.43979e-17 
c_435 M14:DRN B1 2.55268e-17 
c_436 M14:DRN B2 2.10452e-17 
c_437 M14:DRN M9:DRN 2.48382e-18 
c_438 M14:DRN M8:GATE 1.38616e-18 
c_439 M14:DRN M7:DRN 2.32949e-19 
c_440 M14:DRN M7:GATE 1.31418e-19 
c_441 M14:DRN M7:SRC 2.52703e-18 
c_442 M14:DRN M20:SRC 6.57876e-19 
c_443 M14:DRN M11:SRC 9.40805e-19 
c_444 M14:DRN M22:SRC 2.68042e-19 
c_445 M14:DRN M3:DRN 2.56004e-18 
c_446 M14:DRN M14:GATE 1.68073e-17 
c_447 M14:DRN 0 4.18305e-19 
c_448 M6:SRC M10:DRN 6.02021e-18 
c_449 M6:SRC M1:SRC 1.55842e-17 
c_450 M6:SRC M1:DRN 4.26123e-18 
c_451 M6:SRC GND 2.81855e-18 
c_452 M6:SRC M17:SRC 1.66009e-18 
c_453 M6:SRC M1:GATE 5.19446e-19 
c_454 M6:SRC N_4:2 7.87351e-18 
c_455 M6:SRC M10:GATE 4.66634e-19 
c_456 M6:SRC M2:SRC 4.09002e-18 
c_457 M6:SRC A3 9.82188e-17 
c_458 M6:SRC VDD 1.65213e-17 
c_459 M6:SRC M3:GATE 2.09284e-17 
c_460 M6:SRC M4:DRN 3.01936e-18 
c_461 M6:SRC M4:GATE 2.74581e-18 
c_462 M6:SRC M15:GATE 8.7271e-18 
c_463 M6:SRC M5:DRN 2.7132e-18 
c_464 M6:SRC A1 1.83772e-18 
c_465 M6:SRC M5:GATE 9.93674e-18 
c_466 M6:SRC M16:GATE 1.37516e-17 
c_467 M6:SRC M17:DRN 4.73483e-18 
c_468 M6:SRC M17:GATE 5.75474e-19 
c_469 M6:SRC M6:GATE 8.99555e-19 
c_470 M6:SRC B1 1.2376e-17 
c_471 M6:SRC B2 9.00782e-20 
c_472 M6:SRC M2:GATE 4.16059e-19 
c_473 M6:SRC M12:DRN 9.18129e-19 
c_474 M6:SRC M12:SRC 5.13402e-19 
c_475 M6:SRC A2 1.19761e-16 
c_476 M6:SRC 0 9.33879e-20 

.ENDS
