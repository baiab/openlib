
.subckt NR2D1  A1 A2 ZN
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.06318p as=0.12636p l=0.09u nrd=0.217 nrs=0.433 pd=0.774u ps=1.548u sa=5.58e-07 sb=2.34e-07 w=0.54u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.12636p as=0.06318p l=0.09u nrd=0.433 nrs=0.217 pd=1.548u ps=0.774u sa=2.34e-07 sb=5.58e-07 w=0.54u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK pch ad=0.0648p as=0.16848p l=0.09u nrd=0.125 nrs=0.325 pd=0.9u ps=1.908u sa=5.04e-07 sb=2.34e-07 w=0.72u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK pch ad=0.20574p as=0.0648p l=0.09u nrd=0.397 nrs=0.125 pd=2.304u ps=0.9u sa=2.34e-07 sb=5.04e-07 w=0.72u 
R1 M1:DRN GND 18.3253
R2 M2:SRC GND 18.4546
R3 M2:BULK M1:BULK 0.001
R4 M2:BULK GND 4.62531
R5 M4:GATE A1 120.68
R6 M4:GATE M2:GATE 276.316
R7 A1 M2:GATE 100.999
R8 M3:GATE A2 124.687
R9 M3:GATE M1:GATE 275.444
R10 A2 M1:GATE 112.775
R11 M4:SRC ZN 18.5122
R12 ZN M2:DRN 9.19978
R13 M2:DRN M1:SRC 0.001
R14 M4:DRN M3:SRC 0.001
R15 VDD M3:DRN 3.63455
R16 M4:BULK M3:BULK 0.001
R17 M3:BULK M3:DRN 0.001
c_1 M1:DRN 0 3.71834e-18 
c_2 M2:SRC 0 4.98877e-19 
c_3 M2:BULK 0 2.92673e-17 
c_4 GND 0 8.30562e-17 
c_5 M4:GATE 0 2.67427e-17 
c_6 A1 GND 1.2761e-17 
c_7 A1 M1:DRN 3.35812e-20 
c_8 A1 M2:BULK 6.94403e-18 
c_9 A1 M2:SRC 6.58651e-18 
c_10 A1 0 3.76881e-18 
c_11 M2:GATE M2:SRC 2.73441e-17 
c_12 M2:GATE M2:BULK 1.91355e-17 
c_13 M2:GATE GND 1.03182e-17 
c_14 M2:GATE 0 7.67478e-21 
c_15 M3:GATE M4:GATE 2.34979e-17 
c_16 M3:GATE 0 2.29729e-17 
c_17 A2 GND 2.18921e-17 
c_18 A2 M1:DRN 3.43686e-17 
c_19 A2 M2:BULK 6.35139e-18 
c_20 A2 M2:SRC 3.35812e-20 
c_21 A2 A1 7.0972e-18 
c_22 A2 M4:GATE 3.65784e-18 
c_23 A2 0 1.89224e-18 
c_24 M1:GATE M2:BULK 1.91464e-17 
c_25 M1:GATE A1 1.19374e-17 
c_26 M1:GATE M2:GATE 5.23042e-18 
c_27 M1:GATE GND 6.18022e-18 
c_28 M1:GATE 0 2.13254e-18 
c_29 M4:SRC M3:GATE 3.68904e-19 
c_30 M4:SRC M4:GATE 1.69476e-17 
c_31 M4:SRC A1 2.82797e-18 
c_32 M4:SRC M2:SRC 2.68184e-18 
c_33 M4:SRC M2:BULK 3.66468e-20 
c_34 M4:SRC M2:GATE 1.55345e-17 
c_35 M4:SRC 0 4.94421e-18 
c_36 ZN GND 9.13623e-17 
c_37 ZN A2 3.53846e-17 
c_38 ZN M1:DRN 2.13566e-19 
c_39 ZN M1:GATE 1.16891e-17 
c_40 ZN M2:GATE 4.1496e-19 
c_41 ZN M2:BULK 6.99978e-18 
c_42 ZN M2:SRC 1.09866e-18 
c_43 ZN A1 1.17332e-16 
c_44 ZN M4:GATE 1.23065e-17 
c_45 ZN M3:GATE 6.54846e-18 
c_46 ZN 0 2.16822e-17 
c_47 M2:DRN GND 2.85057e-18 
c_48 M2:DRN A2 1.72079e-17 
c_49 M2:DRN M1:DRN 2.36936e-19 
c_50 M2:DRN M1:GATE 1.86877e-17 
c_51 M2:DRN M2:GATE 4.95906e-20 
c_52 M2:DRN M2:BULK 1.06469e-17 
c_53 M2:DRN M2:SRC 2.36936e-19 
c_54 M2:DRN A1 3.48345e-17 
c_55 M2:DRN 0 3.02875e-18 
c_56 M4:DRN ZN 1.42768e-18 
c_57 M4:DRN M2:DRN 3.14238e-18 
c_58 VDD M4:DRN 5.35729e-19 
c_59 VDD M4:SRC 1.74944e-18 
c_60 VDD M3:GATE 1.24579e-17 
c_61 VDD M4:GATE 8.2397e-18 
c_62 VDD ZN 3.43232e-17 
c_63 VDD A2 1.67743e-17 
c_64 VDD A1 1.92808e-18 
c_65 VDD M2:DRN 3.33491e-19 
c_66 VDD 0 7.97141e-17 
c_67 M3:BULK M3:GATE 4.24345e-18 
c_68 M3:BULK M4:GATE 4.57116e-18 
c_69 M3:BULK ZN 1.08781e-17 
c_70 M3:BULK A2 1.08948e-17 
c_71 M3:BULK A1 7.68857e-18 
c_72 M3:DRN M4:DRN 6.53018e-18 
c_73 M3:DRN M4:SRC 1.05143e-17 
c_74 M3:DRN M3:GATE 3.92324e-17 
c_75 M3:DRN M4:GATE 1.23059e-17 
c_76 M3:DRN ZN 1.63271e-18 
c_77 M3:DRN A2 1.6614e-17 
c_78 M3:DRN A1 5.68625e-19 
c_79 M3:DRN M2:DRN 7.14911e-19 
c_80 M3:DRN 0 3.65032e-17 

.ENDS
