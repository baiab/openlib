
.subckt SDFCSND4  SI D SE CP CDN SDN Q QN
MM9 M9:DRN M9:GATE M9:SRC M9:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=1.071e-06 sb=1.413e-06 w=0.54u 
MM10 M10:DRN M10:GATE M10:SRC M10:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=7.47e-07 sb=1.737e-06 w=0.54u 
MM12 M12:DRN M12:GATE M12:SRC M12:BULK nch ad=0.06318p as=0.0972p l=0.09u nrd=0.217 nrs=0.334 pd=0.774u ps=1.764u sa=1.44e-07 sb=2.34e-06 w=0.54u 
MM21 M21:DRN M21:GATE M21:SRC M21:BULK nch ad=0.0972p as=0.06561p l=0.09u nrd=0.334 nrs=0.226 pd=1.764u ps=0.8289u sa=4.761e-07 sb=1.44e-07 w=0.54u 
MM14 M14:DRN M14:GATE M14:SRC M14:BULK nch ad=0.08505p as=0.0405p l=0.09u nrd=0.42 nrs=0.2 pd=0.99u ps=0.63u sa=7.83e-07 sb=8.37e-07 w=0.45u 
MM23 M23:DRN M23:GATE M23:SRC M23:BULK nch ad=0.05589p as=0.06237p l=0.09u nrd=0.767 nrs=0.86 pd=0.954u ps=0.8856u sa=2.07e-07 sb=3.663e-07 w=0.27u 
MM16 M16:DRN M16:GATE M16:SRC M16:BULK nch ad=0.0405p as=0.05832p l=0.09u nrd=0.2 nrs=0.288 pd=0.63u ps=0.8046u sa=4.347e-07 sb=1.107e-06 w=0.45u 
MM25 M25:DRN M25:GATE M25:SRC M25:BULK nch ad=0.02997p as=0.04212p l=0.09u nrd=0.925 nrs=1.29 pd=0.603u ps=0.5904u sa=5.67e-07 sb=1.53e-07 w=0.18u 
MM18 M18:DRN M18:GATE M18:SRC M18:BULK nch ad=0.0405p as=0.09315p l=0.09u nrd=0.2 nrs=0.46 pd=0.63u ps=1.314u sa=1.4715e-06 sb=2.07e-07 w=0.45u 
MM2 M2:DRN M2:GATE M2:SRC M2:BULK nch ad=0.03726p as=0.03564p l=0.09u nrd=0.449 nrs=0.428 pd=0.576u ps=0.6426u sa=7.353e-07 sb=2.826e-07 w=0.288u 
MM27 M27:DRN M27:GATE M27:SRC M27:BULK nch ad=0.0162p as=0.05265p l=0.09u nrd=0.5 nrs=1.634 pd=0.36u ps=0.5895u sa=1.071e-06 sb=1.4589e-06 w=0.18u 
MM4 M4:DRN M4:GATE M4:SRC M4:BULK nch ad=0.0162p as=0.0162p l=0.09u nrd=0.5 nrs=0.5 pd=0.36u ps=0.36u sa=8.01e-07 sb=1.7334e-06 w=0.18u 
MM29 M29:DRN M29:GATE M29:SRC M29:BULK nch ad=0.03078p as=0.10044p l=0.09u nrd=0.263 nrs=0.86 pd=0.522u ps=1.1205u sa=5.859e-07 sb=6.741e-07 w=0.342u 
MM6 M6:DRN M6:GATE M6:SRC M6:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=1.953e-06 sb=5.31e-07 w=0.54u 
MM8 M8:DRN M8:GATE M8:SRC M8:BULK nch ad=0.06318p as=0.06075p l=0.09u nrd=0.217 nrs=0.209 pd=0.774u ps=0.927u sa=1.35e-06 sb=1.134e-06 w=0.54u 
MM11 M11:DRN M11:GATE M11:SRC M11:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=4.68e-07 sb=2.016e-06 w=0.54u 
MM20 M20:DRN M20:GATE M20:SRC M20:BULK nch ad=0.11178p as=0.06723p l=0.09u nrd=0.383 nrs=0.231 pd=1.494u ps=0.945u sa=2.07e-07 sb=5.04e-07 w=0.54u 
MM13 M13:DRN M13:GATE M13:SRC M13:BULK nch ad=0.08505p as=0.0405p l=0.09u nrd=0.42 nrs=0.2 pd=0.99u ps=0.63u sa=1.1853e-06 sb=4.77e-07 w=0.45u 
MM22 M22:DRN M22:GATE M22:SRC M22:BULK nch ad=0.02673p as=0.02997p l=0.09u nrd=0.828 nrs=0.925 pd=0.3897u ps=0.603u sa=1.53e-07 sb=7.92e-07 w=0.18u 
MM15 M15:DRN M15:GATE M15:SRC M15:BULK nch ad=0.0405p as=0.02835p l=0.09u nrd=0.412 nrs=0.286 pd=0.5634u ps=0.495u sa=5.04e-07 sb=1.431e-06 w=0.315u 
MM24 M24:DRN M24:GATE M24:SRC M24:BULK nch ad=0.06966p as=0.05751p l=0.09u nrd=0.318 nrs=0.261 pd=1.0143u ps=0.7191u sa=2.52e-07 sb=4.68e-07 w=0.468u 
MM17 M17:DRN M17:GATE M17:SRC M17:BULK nch ad=0.02835p as=0.11097p l=0.09u nrd=0.286 nrs=1.12 pd=0.495u ps=1.494u sa=2.34e-07 sb=1.701e-06 w=0.315u 
MM1 M1:DRN M1:GATE M1:SRC M1:BULK nch ad=0.03888p as=0.02187p l=0.09u nrd=1.2 nrs=0.685 pd=0.792u ps=0.4014u sa=1.1781e-06 sb=2.16e-07 w=0.18u 
MM26 M26:DRN M26:GATE M26:SRC M26:BULK nch ad=0.09315p as=0.05751p l=0.09u nrd=0.46 nrs=0.286 pd=1.314u ps=0.9774u sa=2.07e-07 sb=2.538e-07 w=0.45u 
MM19 M19:DRN M19:GATE M19:SRC M19:BULK nch ad=0.11178p as=0.06723p l=0.09u nrd=0.383 nrs=0.231 pd=1.494u ps=0.945u sa=5.04e-07 sb=2.07e-07 w=0.54u 
MM3 M3:DRN M3:GATE M3:SRC M3:BULK nch ad=0.04455p as=0.03078p l=0.09u nrd=0.378 nrs=0.263 pd=0.684u ps=0.522u sa=9.405e-07 sb=3.375e-07 w=0.342u 
MM28 M28:DRN M28:GATE M28:SRC M28:BULK nch ad=0.0162p as=0.02349p l=0.09u nrd=0.5 nrs=0.714 pd=0.36u ps=0.3906u sa=5.31e-07 sb=2.0061e-06 w=0.18u 
MM5 M5:DRN M5:GATE M5:SRC M5:BULK nch ad=0.11178p as=0.06318p l=0.09u nrd=0.383 nrs=0.217 pd=1.494u ps=0.774u sa=2.277e-06 sb=2.07e-07 w=0.54u 
MM7 M7:DRN M7:GATE M7:SRC M7:BULK nch ad=0.06075p as=0.06318p l=0.09u nrd=0.209 nrs=0.217 pd=0.927u ps=0.774u sa=1.674e-06 sb=8.1e-07 w=0.54u 
MM51 M51:DRN M51:GATE M51:SRC M51:BULK pch ad=0.07776p as=0.08424p l=0.09u nrd=0.15 nrs=0.162 pd=1.107u ps=0.954u sa=2.8188e-06 sb=8.1e-07 w=0.72u 
MM44 M44:DRN M44:GATE M44:SRC M44:BULK pch ad=0.02187p as=0.03969p l=0.09u nrd=0.3 nrs=0.54 pd=0.432u ps=0.5184u sa=7.83e-07 sb=7.92e-07 w=0.27u 
MM37 M37:DRN M37:GATE M37:SRC M37:BULK pch ad=0.04698p as=0.04455p l=0.09u nrd=0.36 nrs=0.343 pd=0.6984u ps=0.6237u sa=8.1e-07 sb=3.555e-07 w=0.36u 
MM53 M53:DRN M53:GATE M53:SRC M53:BULK pch ad=0.07776p as=0.08424p l=0.09u nrd=0.15 nrs=0.162 pd=1.107u ps=0.954u sa=2.1177e-06 sb=1.413e-06 w=0.72u 
MM46 M46:DRN M46:GATE M46:SRC M46:BULK pch ad=0.14904p as=0.08181p l=0.09u nrd=0.287 nrs=0.158 pd=1.854u ps=1.116u sa=2.07e-07 sb=4.608e-07 w=0.72u 
MM39 M39:DRN M39:GATE M39:SRC M39:BULK pch ad=0.05994p as=0.10449p l=0.09u nrd=0.228 nrs=0.398 pd=0.747u ps=1.062u sa=8.964e-07 sb=3.474e-06 w=0.513u 
MM55 M55:DRN M55:GATE M55:SRC M55:BULK pch ad=0.07776p as=0.08424p l=0.09u nrd=0.15 nrs=0.162 pd=1.107u ps=0.954u sa=1.3176e-06 sb=2.016e-06 w=0.72u 
MM48 M48:DRN M48:GATE M48:SRC M48:BULK pch ad=0.09153p as=0.07695p l=0.09u nrd=0.231 nrs=0.193 pd=1.2096u ps=0.8901u sa=3.105e-07 sb=4.68e-07 w=0.63u 
MM57 M57:DRN M57:GATE M57:SRC M57:BULK pch ad=0.12069p as=0.06723p l=0.09u nrd=0.354 nrs=0.197 pd=1.584u ps=1.017u sa=2.07e-07 sb=6.651e-07 w=0.585u 
MM30 M30:DRN M30:GATE M30:SRC M30:BULK pch ad=0.07452p as=0.04374p l=0.09u nrd=0.575 nrs=0.336 pd=1.134u ps=0.6786u sa=2.07e-07 sb=4.941e-07 w=0.36u 
MM32 M32:DRN M32:GATE M32:SRC M32:BULK pch ad=0.05184p as=0.0324p l=0.09u nrd=0.821 nrs=0.515 pd=0.918u ps=0.4896u sa=1.134e-06 sb=2.07e-07 w=0.252u 
MM41 M41:DRN M41:GATE M41:SRC M41:BULK pch ad=0.05022p as=0.0972p l=0.09u nrd=0.271 nrs=0.52 pd=0.666u ps=1.485u sa=4.68e-07 sb=4.077e-06 w=0.432u 
MM34 M34:DRN M34:GATE M34:SRC M34:BULK pch ad=0.03807p as=0.06642p l=0.09u nrd=0.527 nrs=0.909 pd=0.5985u ps=1.062u sa=5.418e-07 sb=3.627e-07 w=0.27u 
MM50 M50:DRN M50:GATE M50:SRC M50:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=3.1284e-06 sb=5.31e-07 w=0.72u 
MM43 M43:DRN M43:GATE M43:SRC M43:BULK pch ad=0.05994p as=0.11259p l=0.09u nrd=0.228 nrs=0.427 pd=0.747u ps=1.0332u sa=1.6596e-06 sb=2.754e-06 w=0.513u 
MM36 M36:DRN M36:GATE M36:SRC M36:BULK pch ad=0.06156p as=0.10854p l=0.09u nrd=0.261 nrs=0.46 pd=0.9846u ps=1.746u sa=1.611e-07 sb=2.655e-07 w=0.486u 
MM52 M52:DRN M52:GATE M52:SRC M52:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=2.4489e-06 sb=1.134e-06 w=0.72u 
MM45 M45:DRN M45:GATE M45:SRC M45:BULK pch ad=0.12636p as=0.08181p l=0.09u nrd=0.244 nrs=0.158 pd=1.872u ps=1.116u sa=4.95e-07 sb=1.701e-07 w=0.72u 
MM38 M38:DRN M38:GATE M38:SRC M38:BULK pch ad=0.05994p as=0.10449p l=0.09u nrd=0.228 nrs=0.398 pd=0.747u ps=1.062u sa=1.3239e-06 sb=3.078e-06 w=0.513u 
MM54 M54:DRN M54:GATE M54:SRC M54:BULK pch ad=0.08424p as=0.07776p l=0.09u nrd=0.162 nrs=0.15 pd=0.954u ps=1.107u sa=1.7082e-06 sb=1.737e-06 w=0.72u 
MM47 M47:DRN M47:GATE M47:SRC M47:BULK pch ad=0.12312p as=0.08748p l=0.09u nrd=0.238 nrs=0.169 pd=2.124u ps=1.0179u sa=5.49e-07 sb=1.44e-07 w=0.72u 
MM56 M56:DRN M56:GATE M56:SRC M56:BULK pch ad=0.08424p as=0.15795p l=0.09u nrd=0.162 nrs=0.304 pd=0.954u ps=1.4508u sa=7.731e-07 sb=2.34e-06 w=0.72u 
MM49 M49:DRN M49:GATE M49:SRC M49:BULK pch ad=0.14904p as=0.08424p l=0.09u nrd=0.287 nrs=0.162 pd=1.854u ps=0.954u sa=3.4803e-06 sb=2.07e-07 w=0.72u 
MM58 M58:DRN M58:GATE M58:SRC M58:BULK pch ad=0.06723p as=0.07209p l=0.09u nrd=0.197 nrs=0.211 pd=1.017u ps=1.0143u sa=4.86e-07 sb=3.069e-07 w=0.585u 
MM31 M31:DRN M31:GATE M31:SRC M31:BULK pch ad=0.0324p as=0.02187p l=0.09u nrd=0.448 nrs=0.3 pd=0.5094u ps=0.432u sa=5.31e-07 sb=1.044e-06 w=0.27u 
MM40 M40:DRN M40:GATE M40:SRC M40:BULK pch ad=0.05994p as=0.11502p l=0.09u nrd=0.228 nrs=0.438 pd=0.747u ps=1.764u sa=4.815e-07 sb=3.798e-06 w=0.513u 
MM33 M33:DRN M33:GATE M33:SRC M33:BULK pch ad=0.0324p as=0.02835p l=0.09u nrd=0.633 nrs=0.564 pd=0.4995u ps=0.4554u sa=4.797e-07 sb=8.55e-07 w=0.225u 
MM42 M42:DRN M42:GATE M42:SRC M42:BULK pch ad=0.05022p as=0.0972p l=0.09u nrd=0.271 nrs=0.52 pd=0.666u ps=1.485u sa=1.44e-07 sb=4.401e-06 w=0.432u 
MM35 M35:DRN M35:GATE M35:SRC M35:BULK pch ad=0.05589p as=0.06642p l=0.09u nrd=0.767 nrs=0.909 pd=0.954u ps=1.062u sa=5.832e-07 sb=2.07e-07 w=0.27u 
R1 M25:DRN M22:SRC 4.04798e-10
R2 M44:DRN M31:SRC 0.001
R3 M44:GATE M30:DRN 215.613
R4 M44:GATE M24:GATE 325.97
R5 M44:GATE M23:DRN 207.954
R6 M30:DRN M24:GATE 272.766
R7 M30:DRN M23:DRN 43.3872
R8 M24:GATE M23:DRN 263.076
R9 M31:GATE M25:GATE 253.121
R10 M31:GATE SI 104.484
R11 SI M25:GATE 59.9446
R12 M48:SRC M24:SRC 36.5158
R13 M48:SRC M47:SRC 0.001
R14 M24:SRC M21:SRC 0.001
R15 M46:GATE M20:GATE 289.061
R16 M46:GATE CP 116.641
R17 CP M20:GATE 97.828
R18 M47:GATE M21:GATE 297.009
R19 M47:GATE D 92.3837
R20 D M21:GATE 75.4797
R21 M48:GATE M30:GATE 217.08
R22 M30:GATE M23:GATE 253.432
R23 M30:GATE SE 93.0152
R24 SE M23:GATE 66.6115
R25 M23:GATE M22:GATE 163.08
R26 M13:SRC M18:DRN 0.001
R27 M14:SRC M16:DRN 0.001
R28 M3:SRC M29:DRN 0.001
R29 M15:SRC M17:DRN 0.001
R30 M27:DRN M4:DRN 0.001
R31 M26:DRN M22:DRN 28.6516
R32 M24:DRN M22:DRN 3.54388e-10
R33 M4:SRC M28:DRN 0.001
R34 M33:DRN M34:DRN 7.6e-10
R35 M34:DRN M35:DRN 36.5127
R36 M33:GATE M45:GATE 287.138
R37 M33:GATE M37:GATE 97.5975
R38 M37:GATE M45:GATE 717.781
R39 M37:GATE M1:GATE 88.4329
R40 M26:GATE M19:GATE 169.56
R41 M45:GATE M19:GATE 226.27
R42 M45:GATE M20:DRN 225.219
R43 M45:GATE M46:DRN 227.86
R44 M46:DRN M19:GATE 186.362
R45 M46:DRN M20:DRN 45.3801
R46 M19:GATE M20:DRN 184.202
R47 M45:DRN M19:DRN 43.845
R48 M45:DRN M36:GATE 170.596
R49 M45:DRN M28:GATE 316.456
R50 M36:GATE M19:DRN 170.074
R51 M36:GATE M28:GATE 314.021
R52 M32:GATE N_18:1 325.877
R53 M32:GATE M2:GATE 617.773
R54 M2:GATE N_18:1 47.8681
R55 M28:GATE M19:DRN 315.486
R56 M28:GATE N_18:1 44.4992
R57 M57:GATE M28:SRC 345.701
R58 M57:GATE M36:DRN 351.148
R59 M57:GATE M29:GATE 220.607
R60 M36:DRN M28:SRC 45.1016
R61 M36:DRN M29:GATE 132.905
R62 M36:DRN M33:SRC 6.57778e-10
R63 M29:GATE M28:SRC 130.843
R64 M28:SRC M26:SRC 0.001
R65 N_73:1 M48:DRN 19.4624
R66 N_73:1 M36:SRC 18
R67 M48:DRN M44:SRC 0.001
R68 SDN:1 M58:GATE 399
R69 SDN:1 M43:GATE 65.28
R70 M58:GATE M3:GATE 117.51
R71 M43:GATE M18:GATE 229.082
R72 M43:GATE SDN 88.3804
R73 SDN M18:GATE 64.8938
R74 QN M10:DRN 9.2371
R75 QN M53:SRC 18.1828
R76 QN M12:DRN 9.29681
R77 QN M55:SRC 18.406
R78 M55:SRC M56:DRN 0.001
R79 M53:SRC M54:DRN 0.001
R80 M12:DRN M10:DRN 703.543
R81 M12:DRN M11:SRC 0.001
R82 M10:DRN M9:SRC 0.001
R83 Q M8:DRN 9.31172
R84 Q M52:DRN 9.40821
R85 Q M6:DRN 9.23691
R86 Q M50:DRN 9.27762
R87 M52:DRN M50:DRN 605.776
R88 M52:DRN M51:SRC 0.001
R89 M50:DRN M49:SRC 0.001
R90 M8:DRN M6:DRN 704.671
R91 M8:DRN M7:SRC 0.001
R92 M6:DRN M5:SRC 0.001
R93 N_62:1 M34:GATE 57.3759
R94 N_62:1 M4:GATE 93.7139
R95 N_62:1 M57:DRN 18.1657
R96 N_62:1 M58:SRC 18.8885
R97 N_62:1 M2:DRN 18.7293
R98 M58:SRC M2:DRN 1608.05
R99 M58:SRC M37:SRC 2.68658e-10
R100 M34:GATE M4:GATE 196.001
R101 M3:DRN M2:DRN 2.95698e-10
R102 CDN:1 M15:GATE 60.3062
R103 CDN:1 M16:GATE 50.0727
R104 CDN:1 M40:GATE 55.68
R105 CDN:1 M41:GATE 103.277
R106 CDN:1 CDN 24.1852
R107 M35:GATE M27:GATE 94.5
R108 M41:GATE M15:GATE 246.499
R109 M41:GATE CDN 278.381
R110 M27:GATE CDN:2 68.04
R111 CDN M15:GATE 162.554
R112 M15:GATE CDN:2 338.64
R113 GND:1 GND:3 0.592545
R114 GND:1 M21:DRN 1.54168
R115 GND:1 GND:2 0.53703
R116 GND:1 M13:DRN 18
R117 GND:1 M17:SRC 18.4649
R118 GND:2 M25:SRC 18.7538
R119 GND:2 M21:DRN 1.37818
R120 GND:2 GND 0.781066
R121 GND:2 M29:SRC 18.2931
R122 M7:DRN M6:SRC 0.001
R123 M7:DRN M21:DRN 1.42857e-09
R124 M11:DRN M10:SRC 0.001
R125 M11:DRN M21:DRN 1.42857e-09
R126 M12:SRC M21:DRN 1.875e-09
R127 M9:DRN M8:SRC 0.001
R128 M9:DRN M21:DRN 1.42857e-09
R129 M29:BULK M21:DRN 5.26862e-06
R130 M29:BULK M9:BULK 0.001
R131 M29:BULK M23:BULK 0.001
R132 M29:BULK M25:BULK 0.001
R133 M29:BULK M22:BULK 0.001
R134 M29:BULK M24:BULK 0.001
R135 M29:BULK M21:BULK 0.001
R136 M29:BULK M20:BULK 0.001
R137 M29:BULK M19:BULK 0.001
R138 M29:BULK M10:BULK 0.001
R139 M29:BULK M26:BULK 0.001
R140 M29:BULK M28:BULK 0.001
R141 M29:BULK M4:BULK 0.001
R142 M29:BULK M27:BULK 0.001
R143 M29:BULK M3:BULK 0.001
R144 M29:BULK M2:BULK 0.001
R145 M29:BULK M1:BULK 0.001
R146 M29:BULK M17:BULK 0.001
R147 M29:BULK M15:BULK 0.001
R148 M29:BULK M16:BULK 0.001
R149 M29:BULK M14:BULK 0.001
R150 M29:BULK M13:BULK 0.001
R151 M29:BULK M18:BULK 0.001
R152 M29:BULK M12:BULK 0.001
R153 M29:BULK M11:BULK 0.001
R154 M29:BULK M8:BULK 0.001
R155 M29:BULK M7:BULK 0.001
R156 M29:BULK M6:BULK 0.001
R157 M29:BULK M5:BULK 0.001
R158 GND:3 M21:DRN 2.58369
R159 GND:3 M5:DRN 9.28955
R160 M29:SRC M27:SRC 0.001
R161 M13:DRN M21:DRN 5.29952e-10
R162 M13:DRN M14:DRN 0.001
R163 M21:DRN M19:SRC 6.48291e-10
R164 M21:DRN GND 2.27921
R165 M19:SRC M20:SRC 0.001
R166 M25:SRC M23:SRC 0.001
R167 N_56:1 M2:SRC 20.39
R168 N_56:1 M32:SRC 19.8539
R169 N_56:1 M17:GATE 62.7763
R170 N_56:1 M14:GATE 75.0416
R171 N_56:1 M39:GATE 81.5638
R172 N_56:1 M42:GATE 75.4606
R173 M39:GATE M14:GATE 224.211
R174 M42:GATE M17:GATE 174.638
R175 M32:SRC M2:SRC 390.735
R176 M32:SRC M37:DRN 0.001
R177 M2:SRC M1:SRC 8.22222e-10
R178 N_15:1 N_15:3 16.8524
R179 N_15:1 M8:GATE 49.4463
R180 N_15:1 M7:GATE 137.142
R181 N_15:1 N_15:2 31.4452
R182 N_15:1 M52:GATE 66.96
R183 N_15:1 M51:GATE 163.515
R184 N_15:2 M7:GATE 135.203
R185 N_15:2 M6:GATE 56.16
R186 N_15:2 M5:GATE 83.6558
R187 N_15:2 M51:GATE 161.204
R188 N_15:2 M50:GATE 66.96
R189 N_15:2 M49:GATE 99.7434
R190 N_15:3 M41:DRN 18.9343
R191 N_15:3 M15:DRN 19.263
R192 N_15:3 M39:DRN 18.5214
R193 N_15:3 M13:GATE 71.4006
R194 N_15:3 M38:GATE 85.1383
R195 M51:GATE M7:GATE 703.056
R196 M49:GATE M5:GATE 374.592
R197 M39:DRN M41:DRN 1293.07
R198 M39:DRN M40:DRN 0.001
R199 M38:GATE M15:DRN 5371.01
R200 M38:GATE M13:GATE 231.077
R201 M41:DRN M42:DRN 0.001
R202 M13:GATE M15:DRN 4504.36
R203 M15:DRN M16:SRC 1.94241e-10
R204 N_13:1 M1:DRN 24.1229
R205 N_13:1 M32:DRN 24.7104
R206 N_13:1 M18:SRC 19.8327
R207 N_13:1 M43:DRN 18.5613
R208 N_13:1 N_13:2 15.1609
R209 N_13:2 N_13:3 32.0357
R210 N_13:2 M12:GATE 50.3082
R211 N_13:2 M11:GATE 139.717
R212 N_13:2 M56:GATE 66.96
R213 N_13:2 M55:GATE 166.586
R214 N_13:3 M9:GATE 83.6558
R215 N_13:3 M10:GATE 56.16
R216 N_13:3 M11:GATE 133.497
R217 N_13:3 M54:GATE 66.96
R218 N_13:3 M53:GATE 99.7434
R219 N_13:3 M55:GATE 159.169
R220 M55:GATE M11:GATE 694.183
R221 M53:GATE M9:GATE 374.592
R222 M43:DRN M38:DRN 0.001
R223 M18:SRC M1:DRN 621.875
R224 M18:SRC M32:DRN 637.02
R225 M32:DRN M1:DRN 164.195
R226 VDD:1 M47:DRN 45.2949
R227 VDD:1 VDD:3 0.345641
R228 VDD:1 M57:SRC 2.35432
R229 VDD:1 M42:SRC 18.1708
R230 VDD:1 VDD:2 0.360114
R231 VDD:2 M57:SRC 1.33145
R232 VDD:2 M38:SRC 18.2899
R233 VDD:2 M56:SRC 18.2567
R234 VDD:2 M49:DRN 10.7909
R235 VDD:3 M47:DRN 1.93716
R236 VDD:3 M31:DRN 18.7088
R237 VDD:3 VDD 0.704189
R238 VDD:3 M35:SRC 18
R239 VDD:3 M57:SRC 11.2379
R240 M58:BULK M47:DRN 5.2446e-06
R241 M58:BULK M46:SRC 0.00514403
R242 M58:BULK M53:DRN 0.00561167
R243 M58:BULK M35:SRC 0.00237417
R244 M58:BULK M57:SRC 0.00561167
R245 M58:BULK M56:SRC 0.00237417
R246 M58:BULK M55:DRN 0.00561167
R247 M58:BULK M51:DRN 0.00561167
R248 M58:BULK M49:BULK 0.001
R249 M58:BULK M54:BULK 0.001
R250 M58:BULK M30:BULK 0.001
R251 M58:BULK M31:BULK 0.001
R252 M58:BULK M44:BULK 0.001
R253 M58:BULK M53:BULK 0.001
R254 M58:BULK M48:BULK 0.001
R255 M58:BULK M47:BULK 0.001
R256 M58:BULK M46:BULK 0.001
R257 M58:BULK M45:BULK 0.001
R258 M58:BULK M36:BULK 0.001
R259 M58:BULK M33:BULK 0.001
R260 M58:BULK M34:BULK 0.001
R261 M58:BULK M35:BULK 0.001
R262 M58:BULK M57:BULK 0.001
R263 M58:BULK M37:BULK 0.001
R264 M58:BULK M32:BULK 0.001
R265 M58:BULK M42:BULK 0.001
R266 M58:BULK M41:BULK 0.001
R267 M58:BULK M40:BULK 0.001
R268 M58:BULK M39:BULK 0.001
R269 M58:BULK M38:BULK 0.001
R270 M58:BULK M43:BULK 0.001
R271 M58:BULK M56:BULK 0.001
R272 M58:BULK M55:BULK 0.001
R273 M58:BULK M52:BULK 0.001
R274 M58:BULK M51:BULK 0.001
R275 M58:BULK M50:BULK 0.001
R276 VDD M47:DRN 2.38408
R277 M55:DRN M54:SRC 0.001
R278 M55:DRN M57:SRC 6.36364e-10
R279 M53:DRN M52:SRC 0.001
R280 M53:DRN M57:SRC 1.01515e-09
R281 M51:DRN M50:SRC 0.001
R282 M51:DRN M57:SRC 6.16601e-10
R283 M56:SRC M57:SRC 4.61538e-10
R284 M56:SRC M43:SRC 0.001
R285 M49:DRN M57:SRC 80.5802
R286 M57:SRC M47:DRN 1.55e-09
R287 M57:SRC M58:DRN 0.001
R288 M38:SRC M39:SRC 0.001
R289 M42:SRC M40:SRC 1.85859e-09
R290 M40:SRC M41:SRC 0.001
R291 M35:SRC M47:DRN 4.61538e-10
R292 M35:SRC M34:SRC 0.001
R293 M47:DRN M46:SRC 5.83333e-10
R294 M46:SRC M45:SRC 0.001
R295 M31:DRN M30:SRC 0.001
c_1 M25:DRN 0 6.36944e-20 
c_2 M22:SRC 0 5.12627e-20 
c_3 M44:DRN M25:DRN 9.3013e-19 
c_4 M44:DRN M22:SRC 1.48869e-19 
c_5 M44:DRN 0 2.84906e-19 
c_6 M44:GATE 0 4.7343e-18 
c_7 M30:DRN M22:SRC 9.98145e-19 
c_8 M30:DRN 0 2.13076e-19 
c_9 M24:GATE 0 5.30103e-17 
c_10 M23:DRN M25:DRN 3.81485e-18 
c_11 M23:DRN M22:SRC 5.4907e-20 
c_12 M23:DRN 0 5.7166e-20 
c_13 M31:GATE M30:DRN 8.48444e-18 
c_14 M31:GATE M44:GATE 2.04593e-17 
c_15 M31:GATE 0 1.4071e-17 
c_16 SI M25:DRN 1.67676e-19 
c_17 SI M23:DRN 8.06572e-17 
c_18 SI M44:DRN 2.74271e-18 
c_19 SI M44:GATE 4.21641e-18 
c_20 SI 0 1.42163e-17 
c_21 M25:GATE M30:DRN 4.93618e-18 
c_22 M25:GATE M22:SRC 9.12485e-18 
c_23 M25:GATE M23:DRN 1.52522e-19 
c_24 M25:GATE M44:GATE 7.44594e-18 
c_25 M25:GATE 0 1.01742e-18 
c_26 M48:SRC M30:DRN 2.92155e-18 
c_27 M48:SRC M44:GATE 1.06851e-18 
c_28 M48:SRC 0 1.41886e-17 
c_29 M24:SRC M30:DRN 4.29568e-17 
c_30 M24:SRC M24:GATE 2.58356e-17 
c_31 M24:SRC M44:GATE 9.18795e-19 
c_32 M24:SRC 0 1.53275e-17 
c_33 M46:GATE 0 2.20966e-17 
c_34 CP 0 9.14163e-18 
c_35 M20:GATE 0 2.50538e-18 
c_36 M47:GATE M24:SRC 5.23689e-18 
c_37 M47:GATE M44:GATE 1.60914e-19 
c_38 M47:GATE M48:SRC 1.69197e-17 
c_39 M47:GATE CP 8.27605e-18 
c_40 M47:GATE M46:GATE 2.64459e-18 
c_41 M47:GATE 0 2.17261e-17 
c_42 D M24:GATE 7.51912e-18 
c_43 D M24:SRC 2.52743e-17 
c_44 D M44:GATE 1.04471e-17 
c_45 D M48:SRC 8.43317e-17 
c_46 D CP 7.65225e-17 
c_47 D M46:GATE 1.16526e-18 
c_48 D 0 1.1422e-17 
c_49 M21:GATE M24:GATE 3.14755e-18 
c_50 M21:GATE M24:SRC 6.74698e-18 
c_51 M21:GATE M20:GATE 1.31342e-18 
c_52 M21:GATE CP 1.42101e-17 
c_53 M21:GATE 0 2.29291e-18 
c_54 M48:GATE M30:DRN 1.41053e-17 
c_55 M48:GATE M24:SRC 3.4968e-18 
c_56 M48:GATE M44:DRN 4.26422e-18 
c_57 M48:GATE SI 7.38774e-19 
c_58 M48:GATE M31:GATE 7.39818e-18 
c_59 M48:GATE M44:GATE 7.95817e-18 
c_60 M48:GATE M48:SRC 2.37692e-17 
c_61 M48:GATE 0 3.6123e-18 
c_62 M30:GATE M30:DRN 1.67001e-17 
c_63 M30:GATE M24:SRC 4.43815e-18 
c_64 M30:GATE M23:DRN 8.36146e-18 
c_65 M30:GATE SI 2.79353e-18 
c_66 M30:GATE M31:GATE 7.21188e-18 
c_67 M30:GATE M44:GATE 1.77063e-19 
c_68 M30:GATE 0 1.22106e-17 
c_69 SE M30:DRN 1.1177e-16 
c_70 SE M25:GATE 2.83646e-20 
c_71 SE M24:SRC 3.35273e-19 
c_72 SE M23:DRN 1.84197e-19 
c_73 SE SI 7.40865e-17 
c_74 SE M31:GATE 2.18917e-18 
c_75 SE 0 1.28815e-19 
c_76 M23:GATE M25:GATE 1.74347e-18 
c_77 M23:GATE M24:SRC 1.02484e-20 
c_78 M23:GATE M23:DRN 2.57654e-17 
c_79 M23:GATE SI 2.5664e-18 
c_80 M23:GATE M31:GATE 4.3319e-18 
c_81 M23:GATE M44:GATE 4.68995e-19 
c_82 M23:GATE 0 7.69287e-18 
c_83 M22:GATE M30:DRN 1.00563e-17 
c_84 M22:GATE M25:GATE 9.26763e-18 
c_85 M22:GATE M25:DRN 7.6689e-18 
c_86 M22:GATE M22:SRC 9.01604e-18 
c_87 M22:GATE M24:GATE 5.04253e-18 
c_88 M22:GATE M24:SRC 6.9564e-19 
c_89 M22:GATE 0 4.74486e-18 
c_90 M13:SRC 0 4.16809e-19 
c_91 M14:SRC 0 6.11778e-19 
c_92 M3:SRC 0 6.9984e-20 
c_93 M15:SRC 0 4.57615e-20 
c_94 M27:DRN 0 1.44685e-20 
c_95 M26:DRN M22:GATE 3.80364e-18 
c_96 M26:DRN M24:GATE 1.17221e-18 
c_97 M26:DRN M24:SRC 6.28489e-18 
c_98 M26:DRN M44:GATE 2.98504e-17 
c_99 M26:DRN M48:SRC 5.32372e-17 
c_100 M26:DRN M48:GATE 5.50251e-20 
c_101 M26:DRN 0 3.60752e-17 
c_102 M24:DRN M48:GATE 9.62438e-19 
c_103 M24:DRN M23:GATE 2.98675e-19 
c_104 M24:DRN M30:DRN 1.14158e-17 
c_105 M24:DRN M25:DRN 7.03629e-18 
c_106 M24:DRN M22:SRC 1.66882e-18 
c_107 M24:DRN M22:GATE 9.80641e-18 
c_108 M24:DRN 0 2.14514e-18 
c_109 M22:DRN M22:GATE 1.95133e-17 
c_110 M22:DRN M30:DRN 1.72297e-17 
c_111 M22:DRN M24:GATE 2.17073e-18 
c_112 M22:DRN M24:SRC 4.29084e-19 
c_113 M22:DRN M30:GATE 1.50365e-24 
c_114 M22:DRN M48:GATE 3.00837e-20 
c_115 M22:DRN 0 1.09246e-18 
c_116 M4:SRC 0 3.30626e-20 
c_117 M33:DRN M4:SRC 1.75423e-19 
c_118 M33:DRN 0 2.10969e-18 
c_119 M34:DRN M4:SRC 1.87498e-19 
c_120 M34:DRN 0 9.38699e-18 
c_121 M35:DRN 0 2.31065e-18 
c_122 M33:GATE M46:GATE 1.41757e-19 
c_123 M33:GATE M33:DRN 1.52026e-18 
c_124 M33:GATE M34:DRN 1.53378e-17 
c_125 M33:GATE M35:DRN 1.15521e-17 
c_126 M33:GATE 0 5.80716e-18 
c_127 M37:GATE M34:DRN 1.23273e-16 
c_128 M37:GATE 0 3.70438e-17 
c_129 M1:GATE 0 2.72779e-17 
c_130 M26:GATE M20:GATE 2.29317e-19 
c_131 M26:GATE M26:DRN 4.3177e-17 
c_132 M26:GATE 0 3.35132e-19 
c_133 M45:GATE M26:DRN 2.61021e-23 
c_134 M45:GATE M47:GATE 3.44501e-19 
c_135 M45:GATE M46:GATE 1.91992e-17 
c_136 M45:GATE M35:DRN 6.12444e-20 
c_137 M45:GATE 0 1.52446e-17 
c_138 M46:DRN D 2.62014e-19 
c_139 M46:DRN M47:GATE 1.88539e-18 
c_140 M46:DRN CP 1.16464e-16 
c_141 M46:DRN M46:GATE 1.66054e-17 
c_142 M46:DRN 0 5.23019e-19 
c_143 M19:GATE M21:GATE 2.39331e-19 
c_144 M19:GATE M20:GATE 5.26706e-18 
c_145 M19:GATE M26:DRN 2.28906e-17 
c_146 M19:GATE 0 1.59595e-18 
c_147 M20:DRN M22:DRN 7.42865e-17 
c_148 M20:DRN M21:GATE 3.0614e-18 
c_149 M20:DRN D 8.81046e-18 
c_150 M20:DRN M20:GATE 4.08995e-17 
c_151 M20:DRN M26:DRN 5.34654e-18 
c_152 M20:DRN M47:GATE 1.70648e-18 
c_153 M20:DRN CP 3.83467e-17 
c_154 M20:DRN M46:GATE 1.07868e-17 
c_155 M20:DRN 0 1.17763e-17 
c_156 M45:DRN M19:GATE 3.34434e-21 
c_157 M45:DRN M26:DRN 1.41489e-17 
c_158 M45:DRN M20:DRN 9.14183e-18 
c_159 M45:DRN M46:DRN 1.77409e-18 
c_160 M45:DRN M45:GATE 2.88355e-17 
c_161 M45:DRN M33:GATE 5.43079e-18 
c_162 M45:DRN 0 1.39976e-17 
c_163 M36:GATE M22:DRN 6.26667e-17 
c_164 M36:GATE M33:GATE 1.47527e-17 
c_165 M36:GATE 0 5.31482e-18 
c_166 M32:GATE M37:GATE 5.31775e-18 
c_167 M32:GATE M1:GATE 7.54218e-18 
c_168 M32:GATE 0 3.16225e-17 
c_169 M2:GATE M37:GATE 4.75165e-18 
c_170 M2:GATE 0 9.45557e-18 
c_171 M28:GATE M19:GATE 1.82591e-18 
c_172 M28:GATE M26:DRN 5.65391e-19 
c_173 M28:GATE M26:GATE 1.36164e-17 
c_174 M28:GATE 0 3.5455e-17 
c_175 N_18:1 M19:GATE 3.90247e-18 
c_176 N_18:1 M26:DRN 8.07793e-18 
c_177 N_18:1 M4:SRC 5.41676e-18 
c_178 N_18:1 M27:DRN 2.34765e-18 
c_179 N_18:1 M3:SRC 1.41901e-18 
c_180 N_18:1 M33:GATE 9.96644e-20 
c_181 N_18:1 M37:GATE 5.48857e-20 
c_182 N_18:1 M1:GATE 1.70768e-17 
c_183 N_18:1 0 1.78521e-17 
c_184 M19:DRN M22:DRN 1.84442e-17 
c_185 M19:DRN M19:GATE 7.40326e-17 
c_186 M19:DRN M26:DRN 3.42826e-17 
c_187 M19:DRN M20:DRN 1.68236e-17 
c_188 M19:DRN M26:GATE 1.97677e-17 
c_189 M19:DRN M46:DRN 2.72023e-17 
c_190 M19:DRN M45:GATE 4.24658e-17 
c_191 M19:DRN M33:GATE 1.00201e-19 
c_192 M19:DRN 0 1.25958e-18 
c_193 M57:GATE M45:GATE 1.42591e-20 
c_194 M57:GATE M36:GATE 1.50365e-24 
c_195 M57:GATE N_18:1 1.38807e-18 
c_196 M57:GATE M34:DRN 1.81058e-19 
c_197 M57:GATE M35:DRN 3.48227e-19 
c_198 M57:GATE M3:SRC 3.7276e-18 
c_199 M57:GATE M2:GATE 1.60551e-19 
c_200 M57:GATE M33:GATE 7.6294e-18 
c_201 M57:GATE M37:GATE 2.94687e-19 
c_202 M57:GATE 0 1.45471e-17 
c_203 M36:DRN M19:GATE 1.91362e-23 
c_204 M36:DRN M26:DRN 4.55738e-19 
c_205 M36:DRN M26:GATE 1.48936e-18 
c_206 M36:DRN M45:DRN 2.57376e-17 
c_207 M36:DRN M36:GATE 2.97102e-18 
c_208 M36:DRN N_18:1 1.81612e-16 
c_209 M36:DRN M34:DRN 2.35623e-18 
c_210 M36:DRN M35:DRN 3.62843e-19 
c_211 M36:DRN M33:GATE 3.59783e-17 
c_212 M36:DRN 0 7.673e-20 
c_213 M29:GATE N_18:1 2.88985e-18 
c_214 M29:GATE 0 8.81851e-18 
c_215 M28:SRC M22:DRN 3.74137e-17 
c_216 M28:SRC M19:GATE 1.48769e-17 
c_217 M28:SRC M26:DRN 1.68911e-18 
c_218 M28:SRC M26:GATE 9.0138e-18 
c_219 M28:SRC M45:GATE 1.24472e-18 
c_220 M28:SRC M45:DRN 4.62981e-17 
c_221 M28:SRC M19:DRN 4.13155e-20 
c_222 M28:SRC M36:GATE 7.35427e-18 
c_223 M28:SRC M33:DRN 2.60571e-20 
c_224 M28:SRC M28:GATE 6.84148e-17 
c_225 M28:SRC N_18:1 6.19343e-18 
c_226 M28:SRC M34:DRN 1.03763e-18 
c_227 M28:SRC M27:DRN 1.40022e-18 
c_228 M28:SRC M35:DRN 3.84577e-17 
c_229 M28:SRC M3:SRC 5.19985e-22 
c_230 M28:SRC M33:GATE 3.27519e-17 
c_231 M28:SRC 0 1.87053e-17 
c_232 N_73:1 M24:SRC 4.97168e-17 
c_233 N_73:1 D 8.47855e-18 
c_234 N_73:1 M30:GATE 6.24176e-19 
c_235 N_73:1 M44:GATE 2.04762e-17 
c_236 N_73:1 M48:SRC 5.25373e-18 
c_237 N_73:1 M47:GATE 8.65575e-18 
c_238 N_73:1 M46:DRN 8.65207e-17 
c_239 N_73:1 M45:GATE 9.63468e-18 
c_240 N_73:1 M45:DRN 4.08166e-17 
c_241 N_73:1 M48:GATE 1.028e-17 
c_242 N_73:1 M36:GATE 1.69394e-18 
c_243 N_73:1 M28:SRC 2.18734e-17 
c_244 N_73:1 M33:GATE 6.13746e-18 
c_245 N_73:1 0 2.04237e-17 
c_246 M36:SRC M19:GATE 7.51825e-24 
c_247 M36:SRC M45:GATE 4.07676e-19 
c_248 M36:SRC M45:DRN 5.00525e-17 
c_249 M36:SRC M19:DRN 7.37159e-20 
c_250 M36:SRC M36:GATE 1.62954e-17 
c_251 M36:SRC M28:SRC 7.47673e-20 
c_252 M36:SRC M33:GATE 1.55126e-17 
c_253 M36:SRC 0 1.61172e-18 
c_254 M48:DRN M30:DRN 1.08743e-17 
c_255 M48:DRN M24:SRC 1.88746e-18 
c_256 M48:DRN D 3.91775e-19 
c_257 M48:DRN M30:GATE 1.0576e-17 
c_258 M48:DRN M20:DRN 4.85568e-19 
c_259 M48:DRN M44:GATE 3.70588e-17 
c_260 M48:DRN M48:SRC 1.27581e-19 
c_261 M48:DRN M47:GATE 1.41983e-19 
c_262 M48:DRN M48:GATE 2.07517e-17 
c_263 M48:DRN M28:SRC 5.75932e-20 
c_264 M48:DRN 0 7.83608e-18 
c_265 SDN:1 M57:GATE 1.02081e-18 
c_266 SDN:1 0 3.77911e-17 
c_267 M58:GATE M29:GATE 1.57288e-17 
c_268 M58:GATE M57:GATE 2.81365e-17 
c_269 M58:GATE 0 2.1815e-17 
c_270 M43:GATE M57:GATE 3.71171e-22 
c_271 M43:GATE 0 2.4738e-18 
c_272 SDN 0 1.21603e-17 
c_273 M3:GATE M29:GATE 5.49928e-18 
c_274 M3:GATE 0 4.94882e-17 
c_275 M18:GATE 0 1.37496e-17 
c_276 QN 0 3.07293e-17 
c_277 M55:SRC 0 1.34043e-17 
c_278 M53:SRC 0 1.13125e-17 
c_279 M12:DRN 0 3.05408e-18 
c_280 M10:DRN 0 3.59075e-18 
c_281 Q 0 2.64333e-17 
c_282 M52:DRN 0 4.94645e-19 
c_283 M50:DRN 0 5.08915e-18 
c_284 M8:DRN 0 4.10403e-18 
c_285 M6:DRN 0 1.76834e-18 
c_286 N_62:1 M26:GATE 1.4527e-19 
c_287 N_62:1 M45:GATE 4.64216e-20 
c_288 N_62:1 M45:DRN 9.93226e-19 
c_289 N_62:1 M19:DRN 2.52911e-19 
c_290 N_62:1 M36:GATE 3.66214e-19 
c_291 N_62:1 M28:SRC 1.45481e-17 
c_292 N_62:1 M36:DRN 7.9635e-17 
c_293 N_62:1 M33:DRN 6.3755e-18 
c_294 N_62:1 M28:GATE 1.4765e-17 
c_295 N_62:1 N_18:1 8.19257e-17 
c_296 N_62:1 M34:DRN 2.50077e-17 
c_297 N_62:1 M4:SRC 3.48998e-18 
c_298 N_62:1 M27:DRN 2.91204e-19 
c_299 N_62:1 M35:DRN 7.33575e-17 
c_300 N_62:1 M29:GATE 5.52588e-17 
c_301 N_62:1 M57:GATE 2.7222e-17 
c_302 N_62:1 M3:SRC 2.80995e-19 
c_303 N_62:1 M3:GATE 2.23298e-17 
c_304 N_62:1 M58:GATE 5.72657e-18 
c_305 N_62:1 M2:GATE 2.69215e-18 
c_306 N_62:1 M33:GATE 2.95139e-18 
c_307 N_62:1 M37:GATE 1.1473e-16 
c_308 N_62:1 0 1.74013e-18 
c_309 M57:DRN M36:DRN 4.79302e-20 
c_310 M57:DRN M34:DRN 1.23047e-18 
c_311 M57:DRN M35:DRN 1.91012e-17 
c_312 M57:DRN M29:GATE 2.95633e-17 
c_313 M57:DRN M3:SRC 3.56164e-19 
c_314 M57:DRN M58:GATE 1.47635e-19 
c_315 M57:DRN M33:GATE 5.25086e-18 
c_316 M57:DRN 0 4.62875e-19 
c_317 M58:SRC N_18:1 3.94164e-20 
c_318 M58:SRC M57:GATE 1.47635e-19 
c_319 M58:SRC M3:GATE 1.66013e-17 
c_320 M58:SRC SDN:1 1.01311e-17 
c_321 M58:SRC M2:GATE 3.66872e-18 
c_322 M58:SRC M37:GATE 3.98455e-17 
c_323 M58:SRC M32:GATE 3.20549e-19 
c_324 M58:SRC 0 6.47693e-18 
c_325 M34:GATE M36:GATE 4.45428e-20 
c_326 M34:GATE M28:SRC 1.74701e-19 
c_327 M34:GATE M36:DRN 7.12348e-19 
c_328 M34:GATE M34:DRN 1.15201e-17 
c_329 M34:GATE M35:DRN 7.47305e-18 
c_330 M34:GATE M57:GATE 1.02192e-19 
c_331 M34:GATE M58:GATE 5.762e-21 
c_332 M34:GATE M33:GATE 1.27834e-17 
c_333 M34:GATE 0 6.47322e-18 
c_334 M4:GATE M19:GATE 1.52276e-19 
c_335 M4:GATE M28:SRC 1.37326e-18 
c_336 M4:GATE M28:GATE 4.03672e-18 
c_337 M4:GATE N_18:1 1.38201e-17 
c_338 M4:GATE M57:GATE 4.24038e-20 
c_339 M4:GATE 0 2.61302e-17 
c_340 M3:DRN M1:GATE 3.07998e-19 
c_341 M3:DRN M3:GATE 8.00357e-18 
c_342 M3:DRN M29:GATE 8.07083e-19 
c_343 M3:DRN N_18:1 7.35086e-18 
c_344 M3:DRN M19:DRN 3.61697e-21 
c_345 M3:DRN 0 3.06815e-18 
c_346 M2:DRN N_18:1 2.24677e-17 
c_347 M2:DRN M29:GATE 1.60689e-19 
c_348 M2:DRN M3:GATE 2.08716e-17 
c_349 M2:DRN SDN:1 8.48097e-21 
c_350 M2:DRN M58:GATE 3.15647e-19 
c_351 M2:DRN M32:GATE 2.46545e-19 
c_352 M2:DRN M1:GATE 1.17434e-19 
c_353 M2:DRN 0 4.07934e-18 
c_354 CDN:1 N_18:1 3.77696e-19 
c_355 CDN:1 M14:SRC 8.08676e-19 
c_356 CDN:1 M32:GATE 1.81728e-22 
c_357 CDN:1 0 5.68857e-18 
c_358 M40:GATE 0 5.78189e-18 
c_359 M35:GATE M19:DRN 1.33738e-19 
c_360 M35:GATE M36:GATE 1.36362e-20 
c_361 M35:GATE N_18:1 1.62999e-19 
c_362 M35:GATE M34:DRN 1.06341e-19 
c_363 M35:GATE M34:GATE 8.68074e-18 
c_364 M35:GATE M27:DRN 4.4305e-19 
c_365 M35:GATE M35:DRN 2.55625e-17 
c_366 M35:GATE N_62:1 1.15086e-17 
c_367 M35:GATE M57:DRN 6.92805e-18 
c_368 M35:GATE 0 8.49355e-18 
c_369 M41:GATE M32:GATE 4.34103e-20 
c_370 M41:GATE 0 2.43705e-18 
c_371 M27:GATE M19:DRN 5.06649e-20 
c_372 M27:GATE M28:GATE 5.15362e-19 
c_373 M27:GATE N_18:1 6.30186e-18 
c_374 M27:GATE M34:GATE 1.48711e-17 
c_375 M27:GATE M4:GATE 2.75316e-18 
c_376 M27:GATE M35:DRN 5.62793e-21 
c_377 M27:GATE N_62:1 1.11559e-17 
c_378 M27:GATE M57:DRN 4.66645e-19 
c_379 M27:GATE 0 2.43166e-17 
c_380 CDN N_18:1 5.97387e-20 
c_381 CDN M14:SRC 4.65209e-19 
c_382 CDN 0 2.32014e-17 
c_383 M15:GATE N_18:1 1.82143e-19 
c_384 M15:GATE 0 7.23096e-18 
c_385 M16:GATE 0 1.22627e-18 
c_386 CDN:2 M3:DRN 4.68521e-18 
c_387 CDN:2 M19:DRN 6.73978e-20 
c_388 CDN:2 N_18:1 5.29846e-17 
c_389 CDN:2 M4:GATE 6.74662e-18 
c_390 CDN:2 M35:DRN 3.68438e-19 
c_391 CDN:2 N_62:1 6.70286e-19 
c_392 CDN:2 M57:DRN 2.73613e-21 
c_393 CDN:2 M3:SRC 4.85393e-18 
c_394 CDN:2 M58:SRC 2.67907e-22 
c_395 CDN:2 M2:DRN 1.39444e-18 
c_396 CDN:2 M15:SRC 3.53977e-18 
c_397 CDN:2 M32:GATE 1.22064e-21 
c_398 CDN:2 0 1.8932e-17 
c_399 GND:1 CDN:2 2.03375e-19 
c_400 GND:1 QN 3.72584e-20 
c_401 GND:1 N_18:1 2.66752e-20 
c_402 GND:1 M2:GATE 8.65955e-18 
c_403 GND:1 M15:GATE 1.34479e-18 
c_404 GND:1 M16:GATE 9.42884e-19 
c_405 GND:1 M1:GATE 3.08335e-19 
c_406 GND:1 0 4.41286e-17 
c_407 GND:2 M22:GATE 1.94164e-18 
c_408 GND:2 M23:GATE 4.91076e-18 
c_409 GND:2 M25:GATE 2.354e-18 
c_410 GND:2 M22:DRN 8.06887e-20 
c_411 GND:2 M24:GATE 6.25928e-19 
c_412 GND:2 M21:GATE 5.34068e-20 
c_413 GND:2 M20:GATE 2.06882e-19 
c_414 GND:2 M19:GATE 3.1626e-19 
c_415 GND:2 M26:DRN 2.00095e-19 
c_416 GND:2 CDN:2 4.11314e-18 
c_417 GND:2 SE 1.59556e-18 
c_418 GND:2 SI 1.12011e-18 
c_419 GND:2 M20:DRN 1.58274e-20 
c_420 GND:2 M26:GATE 2.1148e-19 
c_421 GND:2 M28:SRC 6.50998e-21 
c_422 GND:2 N_18:1 6.08903e-17 
c_423 GND:2 M29:GATE 6.81899e-19 
c_424 GND:2 0 3.88567e-17 
c_425 M7:DRN Q 7.80063e-18 
c_426 M7:DRN 0 2.37309e-18 
c_427 M11:DRN QN 8.14513e-18 
c_428 M11:DRN 0 2.37309e-18 
c_429 M12:SRC M19:DRN 6.14115e-24 
c_430 M12:SRC M13:SRC 3.61713e-20 
c_431 M12:SRC 0 4.20339e-18 
c_432 M9:DRN QN 6.41234e-20 
c_433 M9:DRN Q 6.41234e-20 
c_434 M9:DRN 0 3.76568e-18 
c_435 M29:BULK M22:GATE 9.34099e-18 
c_436 M29:BULK M23:GATE 3.02116e-17 
c_437 M29:BULK M25:GATE 8.90191e-18 
c_438 M29:BULK M24:GATE 3.8202e-18 
c_439 M29:BULK M24:SRC 5.06811e-18 
c_440 M29:BULK M21:GATE 6.61931e-18 
c_441 M29:BULK D 9.84148e-19 
c_442 M29:BULK M19:GATE 9.99272e-18 
c_443 M29:BULK M26:DRN 1.28025e-17 
c_444 M29:BULK CDN:2 4.63442e-17 
c_445 M29:BULK SE 4.67771e-19 
c_446 M29:BULK SI 1.00647e-18 
c_447 M29:BULK M26:GATE 9.43851e-18 
c_448 M29:BULK M44:GATE 1.15392e-17 
c_449 M29:BULK CP 1.87637e-18 
c_450 M29:BULK M46:GATE 3.09945e-18 
c_451 M29:BULK M45:GATE 6.89892e-18 
c_452 M29:BULK M45:DRN 7.34577e-18 
c_453 M29:BULK QN 5.41083e-18 
c_454 M29:BULK M28:GATE 9.15238e-18 
c_455 M29:BULK N_18:1 3.51562e-17 
c_456 M29:BULK M29:GATE 1.5515e-17 
c_457 M29:BULK M2:GATE 3.12537e-18 
c_458 M29:BULK M15:GATE 5.60852e-18 
c_459 M29:BULK CDN:1 8.27869e-18 
c_460 M29:BULK M16:GATE 2.97839e-18 
c_461 M29:BULK Q 4.07925e-18 
c_462 M29:BULK M37:GATE 4.24362e-18 
c_463 M29:BULK M27:GATE 5.78675e-18 
c_464 M29:BULK M1:GATE 1.37507e-18 
c_465 M29:BULK CDN 3.24798e-18 
c_466 M29:BULK 0 1.53371e-17 
c_467 GND:3 M22:GATE 1.42031e-18 
c_468 GND:3 M23:GATE 2.80695e-17 
c_469 GND:3 M25:GATE 7.20989e-19 
c_470 GND:3 M22:DRN 2.75527e-18 
c_471 GND:3 M24:DRN 1.59554e-20 
c_472 GND:3 M24:GATE 2.23466e-18 
c_473 GND:3 M24:SRC 2.52988e-18 
c_474 GND:3 M21:GATE 3.34317e-18 
c_475 GND:3 D 1.07553e-18 
c_476 GND:3 M20:GATE 3.15597e-18 
c_477 GND:3 M19:GATE 2.18132e-17 
c_478 GND:3 M26:DRN 2.12062e-16 
c_479 GND:3 CDN:2 7.23255e-17 
c_480 GND:3 M23:DRN 3.40401e-17 
c_481 GND:3 SI 3.66765e-19 
c_482 GND:3 M20:DRN 5.57871e-18 
c_483 GND:3 M26:GATE 1.64436e-18 
c_484 GND:3 CP 6.02836e-19 
c_485 GND:3 M19:DRN 1.13344e-18 
c_486 GND:3 M36:GATE 1.61925e-18 
c_487 GND:3 M28:SRC 7.08406e-18 
c_488 GND:3 M10:DRN 2.7956e-18 
c_489 GND:3 QN 9.19609e-17 
c_490 GND:3 M28:GATE 3.28205e-18 
c_491 GND:3 N_18:1 1.77967e-16 
c_492 GND:3 M27:DRN 2.24382e-19 
c_493 GND:3 M29:GATE 8.11107e-19 
c_494 GND:3 M15:GATE 1.8529e-18 
c_495 GND:3 CDN:1 3.18132e-19 
c_496 GND:3 M16:GATE 2.46064e-18 
c_497 GND:3 M14:SRC 3.10964e-19 
c_498 GND:3 M12:DRN 2.4314e-18 
c_499 GND:3 M8:DRN 2.4314e-18 
c_500 GND:3 Q 1.36694e-16 
c_501 GND:3 M6:DRN 1.35716e-18 
c_502 GND:3 M27:GATE 8.02557e-20 
c_503 GND:3 M1:GATE 6.70793e-19 
c_504 GND:3 0 3.30193e-16 
c_505 M5:DRN M6:DRN 1.68344e-18 
c_506 M5:DRN Q 3.79593e-19 
c_507 M5:DRN 0 4.56688e-18 
c_508 M29:SRC M29:GATE 2.65138e-17 
c_509 M29:SRC CDN:2 4.34973e-17 
c_510 M29:SRC M4:SRC 1.44685e-20 
c_511 M29:SRC N_18:1 8.11408e-18 
c_512 M29:SRC M28:SRC 9.20836e-20 
c_513 M29:SRC M26:DRN 6.51036e-21 
c_514 M29:SRC M19:DRN 1.55373e-20 
c_515 M29:SRC 0 4.41587e-18 
c_516 M13:DRN M19:GATE 1.00587e-19 
c_517 M13:DRN CDN:2 1.08206e-18 
c_518 M13:DRN M19:DRN 6.66377e-21 
c_519 M13:DRN M16:GATE 2.4956e-18 
c_520 M13:DRN M12:DRN 5.10186e-22 
c_521 M13:DRN 0 5.10769e-18 
c_522 M17:SRC CDN:2 1.51924e-17 
c_523 M17:SRC M26:GATE 3.46294e-20 
c_524 M17:SRC M19:DRN 2.77163e-20 
c_525 M17:SRC M28:SRC 1.69521e-22 
c_526 M17:SRC N_18:1 6.62052e-20 
c_527 M17:SRC M3:SRC 3.94947e-22 
c_528 M17:SRC M2:GATE 3.18357e-17 
c_529 M17:SRC M15:GATE 3.34481e-18 
c_530 M17:SRC M16:GATE 1.32409e-19 
c_531 M17:SRC M14:SRC 4.56279e-21 
c_532 M17:SRC M32:GATE 1.02642e-17 
c_533 M17:SRC M1:GATE 9.64768e-19 
c_534 M17:SRC 0 3.11311e-18 
c_535 M21:DRN M22:GATE 2.89798e-17 
c_536 M21:DRN M30:DRN 1.09836e-18 
c_537 M21:DRN M23:GATE 4.26808e-17 
c_538 M21:DRN M25:GATE 1.25769e-18 
c_539 M21:DRN M25:DRN 2.36019e-19 
c_540 M21:DRN M22:SRC 4.23428e-18 
c_541 M21:DRN M22:DRN 4.45707e-18 
c_542 M21:DRN M24:DRN 7.55495e-18 
c_543 M21:DRN M24:GATE 6.92792e-18 
c_544 M21:DRN M24:SRC 1.02198e-17 
c_545 M21:DRN M21:GATE 2.60081e-17 
c_546 M21:DRN D 3.78919e-18 
c_547 M21:DRN M20:GATE 1.38542e-17 
c_548 M21:DRN M19:GATE 4.04587e-17 
c_549 M21:DRN M26:DRN 1.35065e-17 
c_550 M21:DRN CDN:2 2.34465e-16 
c_551 M21:DRN M23:DRN 5.37801e-17 
c_552 M21:DRN M30:GATE 5.11241e-23 
c_553 M21:DRN SE 5.4285e-21 
c_554 M21:DRN M20:DRN 3.99378e-17 
c_555 M21:DRN M26:GATE 2.84836e-17 
c_556 M21:DRN M48:SRC 6.24676e-20 
c_557 M21:DRN CP 1.1077e-18 
c_558 M21:DRN M46:DRN 2.00767e-19 
c_559 M21:DRN M19:DRN 6.44342e-18 
c_560 M21:DRN M48:GATE 3.57258e-22 
c_561 M21:DRN M28:SRC 7.58835e-18 
c_562 M21:DRN M10:DRN 8.05621e-18 
c_563 M21:DRN QN 2.85336e-18 
c_564 M21:DRN M53:SRC 4.42193e-20 
c_565 M21:DRN M28:GATE 3.91081e-18 
c_566 M21:DRN N_18:1 1.59257e-17 
c_567 M21:DRN M4:SRC 6.57671e-19 
c_568 M21:DRN M27:DRN 8.80743e-19 
c_569 M21:DRN M35:GATE 9.35104e-20 
c_570 M21:DRN M29:GATE 1.81548e-18 
c_571 M21:DRN M3:SRC 4.41091e-18 
c_572 M21:DRN M15:SRC 3.27054e-18 
c_573 M21:DRN M15:GATE 6.21854e-20 
c_574 M21:DRN CDN:1 9.18359e-20 
c_575 M21:DRN M16:GATE 6.09307e-18 
c_576 M21:DRN M14:SRC 5.94433e-18 
c_577 M21:DRN M13:SRC 6.04396e-18 
c_578 M21:DRN M12:DRN 1.13251e-17 
c_579 M21:DRN M55:SRC 4.42193e-20 
c_580 M21:DRN M8:DRN 1.13251e-17 
c_581 M21:DRN M52:DRN 4.42193e-20 
c_582 M21:DRN Q 2.7858e-18 
c_583 M21:DRN M6:DRN 1.13251e-17 
c_584 M21:DRN M50:DRN 4.42193e-20 
c_585 M21:DRN 0 2.05969e-16 
c_586 M19:SRC CDN:2 8.87021e-20 
c_587 M19:SRC M26:GATE 6.65617e-19 
c_588 M19:SRC M26:DRN 3.10265e-18 
c_589 M19:SRC M19:GATE 1.21085e-17 
c_590 M19:SRC M20:GATE 5.44328e-18 
c_591 M19:SRC M20:DRN 9.51215e-18 
c_592 M19:SRC M22:GATE 7.99824e-20 
c_593 M19:SRC 0 2.36969e-18 
c_594 M25:SRC M22:GATE 1.62762e-17 
c_595 M25:SRC M23:GATE 2.97622e-17 
c_596 M25:SRC M25:GATE 1.47458e-17 
c_597 M25:SRC M22:SRC 8.41512e-18 
c_598 M25:SRC M22:DRN 1.71705e-20 
c_599 M25:SRC M24:DRN 2.85753e-20 
c_600 M25:SRC M24:GATE 1.72481e-19 
c_601 M25:SRC M24:SRC 2.2655e-20 
c_602 M25:SRC M26:DRN 1.62771e-20 
c_603 M25:SRC M23:DRN 4.71511e-18 
c_604 M25:SRC M30:GATE 6.4657e-23 
c_605 M25:SRC SE 1.24147e-18 
c_606 M25:SRC SI 4.49414e-18 
c_607 M25:SRC M31:GATE 6.12473e-22 
c_608 M25:SRC 0 1.1864e-18 
c_609 GND M23:DRN 1.39715e-20 
c_610 GND M26:DRN 5.66815e-18 
c_611 GND 0 6.37972e-17 
c_612 N_56:1 GND:3 2.99536e-18 
c_613 N_56:1 M21:DRN 2.37586e-19 
c_614 N_56:1 CDN:2 9.69911e-20 
c_615 N_56:1 M29:BULK 9.2571e-18 
c_616 N_56:1 N_18:1 2.62095e-17 
c_617 N_56:1 N_62:1 8.45189e-17 
c_618 N_56:1 M58:SRC 1.02548e-18 
c_619 N_56:1 M2:DRN 8.12829e-19 
c_620 N_56:1 M2:GATE 2.31292e-18 
c_621 N_56:1 M15:GATE 1.3301e-18 
c_622 N_56:1 CDN:1 3.80771e-17 
c_623 N_56:1 M16:GATE 8.00872e-18 
c_624 N_56:1 M14:SRC 2.19985e-18 
c_625 N_56:1 GND:1 1.13762e-18 
c_626 N_56:1 M13:DRN 5.36567e-18 
c_627 N_56:1 M37:GATE 2.96842e-17 
c_628 N_56:1 M32:GATE 2.59492e-17 
c_629 N_56:1 M40:GATE 9.15856e-18 
c_630 N_56:1 M1:GATE 1.42618e-17 
c_631 N_56:1 M41:GATE 1.15489e-19 
c_632 N_56:1 CDN 9.44034e-17 
c_633 N_56:1 0 8.43349e-18 
c_634 M39:GATE M40:GATE 8.8618e-18 
c_635 M39:GATE M41:GATE 2.33676e-19 
c_636 M39:GATE CDN 7.02023e-21 
c_637 M39:GATE 0 1.18164e-17 
c_638 M42:GATE N_18:1 2.73311e-18 
c_639 M42:GATE M15:GATE 1.06575e-17 
c_640 M42:GATE CDN:1 2.14056e-19 
c_641 M42:GATE M37:GATE 2.07339e-19 
c_642 M42:GATE M32:GATE 5.15308e-19 
c_643 M42:GATE M40:GATE 1.82492e-19 
c_644 M42:GATE M41:GATE 4.29978e-18 
c_645 M42:GATE CDN 3.07397e-18 
c_646 M42:GATE 0 3.68181e-18 
c_647 M32:SRC M21:DRN 7.29911e-20 
c_648 M32:SRC CDN:2 4.82749e-23 
c_649 M32:SRC N_18:1 1.67326e-20 
c_650 M32:SRC M58:SRC 7.28765e-19 
c_651 M32:SRC M2:DRN 2.70485e-19 
c_652 M32:SRC M37:GATE 7.49427e-18 
c_653 M32:SRC M32:GATE 2.08749e-17 
c_654 M32:SRC M1:GATE 2.83967e-17 
c_655 M32:SRC 0 3.78471e-18 
c_656 M17:GATE GND:3 7.74709e-19 
c_657 M17:GATE M21:DRN 1.77058e-18 
c_658 M17:GATE CDN:2 4.67243e-18 
c_659 M17:GATE M2:GATE 3.97782e-18 
c_660 M17:GATE M15:GATE 1.16254e-17 
c_661 M17:GATE CDN:1 5.59879e-18 
c_662 M17:GATE M16:GATE 4.82907e-21 
c_663 M17:GATE GND:1 1.39562e-18 
c_664 M17:GATE M17:SRC 2.39184e-17 
c_665 M17:GATE CDN 1.02545e-19 
c_666 M14:GATE GND:3 1.90267e-18 
c_667 M14:GATE M21:DRN 6.08877e-18 
c_668 M14:GATE CDN:2 6.25247e-21 
c_669 M14:GATE M29:BULK 3.13199e-18 
c_670 M14:GATE M15:GATE 7.37926e-20 
c_671 M14:GATE M16:GATE 1.10619e-17 
c_672 M14:GATE GND:1 4.73721e-19 
c_673 M14:GATE M13:DRN 1.60721e-17 
c_674 M14:GATE 0 1.70286e-18 
c_675 M2:SRC M21:DRN 5.20082e-19 
c_676 M2:SRC CDN:2 8.40026e-19 
c_677 M2:SRC M19:DRN 1.4991e-23 
c_678 M2:SRC N_18:1 1.6083e-17 
c_679 M2:SRC N_62:1 8.48943e-19 
c_680 M2:SRC M58:SRC 9.15251e-19 
c_681 M2:SRC M2:DRN 8.28328e-19 
c_682 M2:SRC M2:GATE 1.85376e-17 
c_683 M2:SRC M12:SRC 2.65381e-23 
c_684 M2:SRC M33:GATE 2.28537e-20 
c_685 M2:SRC M37:GATE 1.9179e-17 
c_686 M2:SRC M17:SRC 2.07127e-19 
c_687 M2:SRC M1:GATE 1.15853e-17 
c_688 M2:SRC 0 2.83725e-18 
c_689 N_15:1 GND:3 1.14159e-18 
c_690 N_15:1 M21:DRN 3.66042e-19 
c_691 N_15:1 M29:BULK 7.36318e-18 
c_692 N_15:1 M10:DRN 2.95269e-19 
c_693 N_15:1 QN 3.38796e-18 
c_694 N_15:1 M8:DRN 3.96802e-17 
c_695 N_15:1 M52:DRN 1.49115e-17 
c_696 N_15:1 M7:DRN 1.01575e-17 
c_697 N_15:1 Q 7.30001e-17 
c_698 N_15:1 M6:DRN 1.52448e-17 
c_699 N_15:1 M50:DRN 1.47549e-17 
c_700 N_15:1 M43:GATE 8.15453e-21 
c_701 N_15:2 GND:3 7.62038e-18 
c_702 N_15:2 M21:DRN 1.63248e-19 
c_703 N_15:2 M29:BULK 8.24057e-18 
c_704 N_15:2 M10:DRN 4.50956e-20 
c_705 N_15:2 M8:DRN 1.13071e-17 
c_706 N_15:2 Q 3.13175e-17 
c_707 N_15:2 M6:DRN 2.88499e-17 
c_708 N_15:3 GND:3 8.86669e-18 
c_709 N_15:3 M21:DRN 3.17782e-18 
c_710 N_15:3 CDN:2 1.96497e-19 
c_711 N_15:3 M29:BULK 3.56656e-18 
c_712 N_15:3 QN 1.48931e-16 
c_713 N_15:3 M53:SRC 6.97561e-18 
c_714 N_15:3 M9:DRN 3.0159e-18 
c_715 N_15:3 SDN:1 7.07854e-18 
c_716 N_15:3 N_56:1 2.06308e-16 
c_717 N_15:3 M17:GATE 1.62608e-19 
c_718 N_15:3 M15:GATE 8.73211e-18 
c_719 N_15:3 CDN:1 5.59258e-18 
c_720 N_15:3 M16:GATE 1.76698e-18 
c_721 N_15:3 M14:SRC 2.40259e-18 
c_722 N_15:3 M14:GATE 1.5587e-17 
c_723 N_15:3 GND:1 3.17631e-18 
c_724 N_15:3 M13:DRN 1.02478e-17 
c_725 N_15:3 M13:SRC 4.50271e-18 
c_726 N_15:3 SDN 4.62889e-17 
c_727 N_15:3 M55:SRC 6.13035e-18 
c_728 N_15:3 M8:DRN 1.27849e-18 
c_729 N_15:3 M52:DRN 1.89434e-18 
c_730 N_15:3 Q 8.29081e-17 
c_731 N_15:3 M40:GATE 8.05874e-18 
c_732 N_15:3 M39:GATE 2.87333e-17 
c_733 N_15:3 M41:GATE 4.99493e-18 
c_734 N_15:3 CDN 6.14024e-17 
c_735 N_15:3 M43:GATE 6.62056e-19 
c_736 N_15:3 M42:GATE 2.65124e-18 
c_737 M52:GATE M53:SRC 3.24889e-19 
c_738 M52:GATE M52:DRN 3.37017e-17 
c_739 M52:GATE Q 8.37068e-18 
c_740 M52:GATE 0 3.34592e-18 
c_741 M51:GATE M52:DRN 3.32176e-17 
c_742 M51:GATE Q 1.91505e-17 
c_743 M51:GATE M50:DRN 2.95269e-19 
c_744 M51:GATE 0 1.61199e-18 
c_745 M50:GATE M52:DRN 2.95269e-19 
c_746 M50:GATE Q 2.09068e-17 
c_747 M50:GATE M50:DRN 3.32599e-17 
c_748 M50:GATE 0 1.38525e-18 
c_749 M49:GATE Q 1.13421e-17 
c_750 M49:GATE M6:DRN 8.43608e-18 
c_751 M49:GATE M50:DRN 3.33865e-17 
c_752 M49:GATE M5:DRN 1.89621e-19 
c_753 M49:GATE 0 9.05709e-19 
c_754 M5:GATE M29:BULK 9.62328e-18 
c_755 M5:GATE GND:3 5.32469e-18 
c_756 M5:GATE M6:DRN 1.01227e-17 
c_757 M5:GATE M5:DRN 3.30939e-17 
c_758 M5:GATE M21:DRN 1.12087e-17 
c_759 M6:GATE M29:BULK 4.37323e-18 
c_760 M6:GATE Q 9.81538e-19 
c_761 M6:GATE GND:3 4.68386e-18 
c_762 M6:GATE M6:DRN 2.02974e-17 
c_763 M6:GATE M5:DRN 4.16913e-20 
c_764 M6:GATE M21:DRN 1.94243e-17 
c_765 M6:GATE 0 1.56632e-19 
c_766 M8:GATE M29:BULK 4.6259e-18 
c_767 M8:GATE Q 2.42331e-19 
c_768 M8:GATE GND:3 3.43575e-18 
c_769 M8:GATE M8:DRN 1.59552e-17 
c_770 M8:GATE M21:DRN 2.05768e-17 
c_771 M8:GATE 0 3.38514e-18 
c_772 M7:GATE Q 5.27308e-18 
c_773 M7:GATE M29:BULK 5.71856e-18 
c_774 M7:GATE GND:3 3.14404e-18 
c_775 M7:GATE M8:DRN 1.85454e-17 
c_776 M7:GATE M6:DRN 6.80165e-19 
c_777 M7:GATE M21:DRN 2.09991e-17 
c_778 M39:DRN M21:DRN 5.26306e-19 
c_779 M39:DRN SDN:1 7.63474e-18 
c_780 M39:DRN N_56:1 5.65094e-18 
c_781 M39:DRN M14:SRC 3.45603e-18 
c_782 M39:DRN M14:GATE 7.92188e-18 
c_783 M39:DRN Q 2.96235e-18 
c_784 M39:DRN M40:GATE 1.67484e-17 
c_785 M39:DRN M39:GATE 1.67655e-17 
c_786 M39:DRN M41:GATE 1.47635e-19 
c_787 M39:DRN CDN 4.34074e-19 
c_788 M39:DRN 0 1.17334e-18 
c_789 M38:GATE SDN:1 4.69718e-18 
c_790 M38:GATE N_56:1 5.95552e-19 
c_791 M38:GATE SDN 1.12186e-17 
c_792 M38:GATE M40:GATE 8.73742e-20 
c_793 M38:GATE M39:GATE 4.53133e-18 
c_794 M38:GATE M43:GATE 4.17912e-18 
c_795 M38:GATE 0 2.0659e-18 
c_796 M41:DRN M21:DRN 7.41317e-20 
c_797 M41:DRN CDN:2 2.43108e-18 
c_798 M41:DRN SDN:1 4.12099e-18 
c_799 M41:DRN M32:SRC 3.63979e-21 
c_800 M41:DRN N_56:1 5.93839e-18 
c_801 M41:DRN M15:SRC 5.35535e-18 
c_802 M41:DRN Q 1.33012e-18 
c_803 M41:DRN M40:GATE 1.47635e-19 
c_804 M41:DRN M41:GATE 1.43863e-17 
c_805 M41:DRN CDN 7.20175e-18 
c_806 M41:DRN M42:GATE 1.67814e-17 
c_807 M41:DRN 0 1.14932e-20 
c_808 M13:GATE GND:3 2.09421e-18 
c_809 M13:GATE M21:DRN 6.31176e-18 
c_810 M13:GATE M29:BULK 1.4757e-18 
c_811 M13:GATE M16:GATE 3.5995e-20 
c_812 M13:GATE M14:GATE 7.93607e-19 
c_813 M13:GATE GND:1 5.31032e-19 
c_814 M13:GATE M13:DRN 1.65601e-17 
c_815 M13:GATE M18:GATE 6.16841e-18 
c_816 M13:GATE SDN 2.33474e-17 
c_817 M13:GATE M12:SRC 2.02097e-19 
c_818 M15:DRN GND:3 1.50582e-18 
c_819 M15:DRN M21:DRN 1.68055e-18 
c_820 M15:DRN CDN:2 2.27164e-19 
c_821 M15:DRN QN 9.73105e-20 
c_822 M15:DRN SDN:1 8.6155e-22 
c_823 M15:DRN N_56:1 3.25884e-19 
c_824 M15:DRN M17:GATE 1.60689e-19 
c_825 M15:DRN M15:GATE 1.7373e-17 
c_826 M15:DRN CDN:1 1.22113e-17 
c_827 M15:DRN M16:GATE 4.56527e-18 
c_828 M15:DRN M55:SRC 1.45561e-20 
c_829 M15:DRN CDN 8.8883e-18 
c_830 M15:DRN 0 9.12432e-18 
c_831 M16:SRC M21:DRN 7.11996e-18 
c_832 M16:SRC CDN:2 1.20972e-18 
c_833 M16:SRC M17:GATE 1.78007e-18 
c_834 M16:SRC M15:GATE 3.00392e-18 
c_835 M16:SRC M13:DRN 3.61713e-20 
c_836 M16:SRC M29:SRC 2.10158e-22 
c_837 M16:SRC M17:SRC 1.24385e-18 
c_838 M16:SRC M41:GATE 7.64418e-18 
c_839 M16:SRC 0 4.27612e-23 
c_840 N_13:1 GND:3 1.60524e-16 
c_841 N_13:1 M21:DRN 5.68536e-17 
c_842 N_13:1 GND:2 2.56277e-20 
c_843 N_13:1 M29:BULK 1.02453e-17 
c_844 N_13:1 QN 1.00108e-16 
c_845 N_13:1 N_18:1 3.72268e-19 
c_846 N_13:1 SDN:1 9.63514e-20 
c_847 N_13:1 M2:GATE 1.64595e-17 
c_848 N_13:1 M2:SRC 1.6635e-17 
c_849 N_13:1 M32:SRC 1.84418e-17 
c_850 N_13:1 N_56:1 1.84369e-16 
c_851 N_13:1 M17:GATE 1.94888e-18 
c_852 N_13:1 N_15:3 1.6882e-16 
c_853 N_13:1 M15:SRC 3.1413e-18 
c_854 N_13:1 M41:DRN 4.21954e-19 
c_855 N_13:1 M15:DRN 5.50769e-18 
c_856 N_13:1 M16:SRC 2.14903e-18 
c_857 N_13:1 M14:SRC 2.70876e-18 
c_858 N_13:1 M14:GATE 2.51266e-19 
c_859 N_13:1 M13:DRN 5.88339e-18 
c_860 N_13:1 M13:GATE 6.13904e-18 
c_861 N_13:1 M13:SRC 2.0396e-18 
c_862 N_13:1 M18:GATE 2.66073e-18 
c_863 N_13:1 SDN 7.67041e-17 
c_864 N_13:1 M12:SRC 4.90395e-19 
c_865 N_13:1 M12:DRN 1.89263e-18 
c_866 N_13:1 M55:SRC 1.52777e-18 
c_867 N_13:1 M32:GATE 9.05445e-18 
c_868 N_13:1 M39:GATE 7.76298e-21 
c_869 N_13:1 M38:GATE 1.19239e-17 
c_870 N_13:1 M17:SRC 4.97316e-18 
c_871 N_13:1 M43:GATE 1.17109e-17 
c_872 N_13:1 M42:GATE 1.9162e-18 
c_873 N_13:1 0 4.88631e-17 
c_874 N_13:2 GND:3 1.14159e-18 
c_875 N_13:2 M21:DRN 3.8048e-19 
c_876 N_13:2 M29:BULK 5.68498e-18 
c_877 N_13:2 M10:DRN 1.53543e-17 
c_878 N_13:2 QN 5.58377e-17 
c_879 N_13:2 M53:SRC 1.4766e-17 
c_880 N_13:2 N_15:3 7.45066e-18 
c_881 N_13:2 M13:GATE 8.51507e-20 
c_882 N_13:2 M18:GATE 3.67107e-18 
c_883 N_13:2 SDN 8.34262e-18 
c_884 N_13:2 M12:DRN 3.84525e-17 
c_885 N_13:2 M55:SRC 1.47951e-17 
c_886 N_13:2 M11:DRN 1.01575e-17 
c_887 N_13:2 N_15:1 9.92028e-18 
c_888 N_13:2 M38:GATE 2.25702e-19 
c_889 N_13:2 0 1.44131e-19 
c_890 N_13:3 GND:3 1.56466e-18 
c_891 N_13:3 M21:DRN 5.44161e-20 
c_892 N_13:3 M29:BULK 5.30735e-18 
c_893 N_13:3 M10:DRN 5.89363e-17 
c_894 N_13:3 QN 5.50732e-18 
c_895 N_13:3 N_15:3 6.257e-19 
c_896 N_13:3 M18:GATE 1.05046e-20 
c_897 N_13:3 M12:DRN 9.92363e-18 
c_898 N_13:3 N_15:1 3.54627e-19 
c_899 N_13:3 N_15:2 1.22449e-19 
c_900 N_13:3 M43:GATE 1.22725e-19 
c_901 M56:GATE QN 4.88257e-18 
c_902 M56:GATE SDN:1 5.05843e-19 
c_903 M56:GATE N_15:3 8.85463e-18 
c_904 M56:GATE M18:GATE 3.16311e-18 
c_905 M56:GATE M55:SRC 1.79073e-17 
c_906 M56:GATE M38:GATE 8.21532e-20 
c_907 M56:GATE M43:GATE 1.31009e-18 
c_908 M56:GATE 0 9.68831e-19 
c_909 M55:GATE QN 7.07143e-18 
c_910 M55:GATE M53:SRC 1.47635e-19 
c_911 M55:GATE SDN:1 3.26996e-20 
c_912 M55:GATE N_15:3 1.35819e-19 
c_913 M55:GATE M41:DRN 8.49042e-18 
c_914 M55:GATE M15:DRN 1.46949e-20 
c_915 M55:GATE M12:DRN 3.01843e-18 
c_916 M55:GATE M55:SRC 1.6633e-17 
c_917 M55:GATE M43:GATE 1.88444e-19 
c_918 M55:GATE 0 4.56844e-19 
c_919 M54:GATE QN 8.51889e-18 
c_920 M54:GATE M53:SRC 1.66335e-17 
c_921 M54:GATE N_15:3 9.00898e-18 
c_922 M54:GATE M55:SRC 1.47635e-19 
c_923 M54:GATE M52:GATE 3.15219e-19 
c_924 M54:GATE 0 1.57328e-18 
c_925 M53:GATE QN 3.71403e-18 
c_926 M53:GATE M53:SRC 1.67605e-17 
c_927 M53:GATE N_15:3 1.33461e-17 
c_928 M53:GATE N_15:1 3.77255e-18 
c_929 M53:GATE N_15:2 1.02822e-19 
c_930 M53:GATE M52:GATE 1.86636e-17 
c_931 M53:GATE M51:GATE 1.52009e-19 
c_932 M53:GATE 0 1.65746e-18 
c_933 M43:DRN GND:3 2.02877e-19 
c_934 M43:DRN M21:DRN 4.1345e-19 
c_935 M43:DRN M29:BULK 2.87226e-21 
c_936 M43:DRN SDN:1 8.25246e-18 
c_937 M43:DRN N_15:3 6.74226e-18 
c_938 M43:DRN M39:DRN 4.12353e-20 
c_939 M43:DRN M13:SRC 1.68211e-18 
c_940 M43:DRN SDN 8.76478e-18 
c_941 M43:DRN M55:SRC 4.12353e-20 
c_942 M43:DRN M39:GATE 5.85036e-20 
c_943 M43:DRN M38:GATE 1.67952e-17 
c_944 M43:DRN M43:GATE 1.6671e-17 
c_945 M43:DRN 0 5.06395e-18 
c_946 M11:GATE GND:3 3.14404e-18 
c_947 M11:GATE M21:DRN 2.0952e-17 
c_948 M11:GATE M29:BULK 5.27961e-18 
c_949 M11:GATE QN 2.3561e-18 
c_950 M11:GATE GND:1 6.55561e-20 
c_951 M11:GATE M13:DRN 1.82015e-20 
c_952 M11:GATE M18:GATE 7.23354e-20 
c_953 M11:GATE M12:DRN 2.23796e-17 
c_954 M12:GATE GND:1 2.2835e-20 
c_955 M12:GATE M29:BULK 2.62745e-18 
c_956 M12:GATE QN 1.12304e-18 
c_957 M12:GATE GND:3 3.2197e-18 
c_958 M12:GATE M12:DRN 1.285e-17 
c_959 M12:GATE M13:GATE 7.94157e-20 
c_960 M12:GATE M18:GATE 8.10179e-19 
c_961 M12:GATE M13:DRN 4.2402e-19 
c_962 M12:GATE M21:DRN 2.6274e-17 
c_963 M12:GATE 0 2.49427e-18 
c_964 M10:GATE N_15:1 3.60853e-20 
c_965 M10:GATE M29:BULK 5.28406e-18 
c_966 M10:GATE QN 1.5669e-17 
c_967 M10:GATE M8:GATE 3.89664e-19 
c_968 M10:GATE GND:3 3.14404e-18 
c_969 M10:GATE M12:DRN 2.95269e-19 
c_970 M10:GATE M10:DRN 4.88115e-18 
c_971 M10:GATE M21:DRN 2.10535e-17 
c_972 M10:GATE 0 4.0602e-19 
c_973 M9:GATE GND:3 3.43575e-18 
c_974 M9:GATE M21:DRN 2.06167e-17 
c_975 M9:GATE M29:BULK 6.44984e-18 
c_976 M9:GATE M10:DRN 5.92511e-18 
c_977 M9:GATE QN 7.34917e-18 
c_978 M9:GATE N_15:1 1.48519e-17 
c_979 M9:GATE M8:GATE 4.53526e-18 
c_980 M9:GATE M7:GATE 3.89664e-19 
c_981 M9:GATE 0 2.01811e-18 
c_982 M18:SRC GND:3 2.85383e-18 
c_983 M18:SRC M21:DRN 9.95348e-18 
c_984 M18:SRC QN 2.90602e-20 
c_985 M18:SRC GND:1 1.14752e-19 
c_986 M18:SRC M13:DRN 5.74193e-19 
c_987 M18:SRC M13:GATE 3.46534e-19 
c_988 M18:SRC M18:GATE 3.16986e-17 
c_989 M18:SRC SDN 2.92953e-17 
c_990 M18:SRC M12:SRC 2.45951e-17 
c_991 M18:SRC M12:DRN 9.59572e-20 
c_992 M32:DRN M21:DRN 8.49102e-20 
c_993 M32:DRN QN 1.93556e-17 
c_994 M32:DRN N_18:1 1.89648e-18 
c_995 M32:DRN SDN:1 3.05841e-18 
c_996 M32:DRN M32:SRC 4.36061e-19 
c_997 M32:DRN N_56:1 3.45566e-18 
c_998 M32:DRN N_15:3 5.36684e-17 
c_999 M32:DRN M41:DRN 4.64286e-20 
c_1000 M32:DRN SDN 4.33343e-21 
c_1001 M32:DRN M32:GATE 3.27961e-17 
c_1002 M32:DRN M17:SRC 3.7003e-20 
c_1003 M32:DRN M42:GATE 1.83794e-18 
c_1004 M32:DRN 0 8.8893e-18 
c_1005 M1:DRN M21:DRN 1.79304e-19 
c_1006 M1:DRN SDN:1 1.4771e-20 
c_1007 M1:DRN M2:GATE 2.71045e-17 
c_1008 M1:DRN M2:SRC 4.10645e-19 
c_1009 M1:DRN M32:SRC 9.53016e-19 
c_1010 M1:DRN N_56:1 2.39822e-18 
c_1011 M1:DRN N_15:3 1.04713e-17 
c_1012 M1:DRN M15:SRC 9.40453e-21 
c_1013 M1:DRN GND:1 5.00035e-17 
c_1014 M1:DRN SDN 1.43126e-17 
c_1015 M1:DRN M12:SRC 2.22657e-18 
c_1016 M1:DRN M12:DRN 3.07417e-20 
c_1017 M1:DRN M32:GATE 5.00756e-18 
c_1018 M1:DRN M17:SRC 4.32793e-18 
c_1019 M1:DRN 0 2.39552e-17 
c_1020 VDD:1 M58:GATE 7.07529e-21 
c_1021 VDD:1 M32:DRN 7.94223e-19 
c_1022 VDD:1 N_56:1 5.11532e-17 
c_1023 VDD:1 N_15:3 1.35343e-18 
c_1024 VDD:1 SDN 5.94871e-21 
c_1025 VDD:1 N_13:1 8.01809e-19 
c_1026 VDD:1 Q 1.18707e-19 
c_1027 VDD:1 M37:GATE 1.41607e-18 
c_1028 VDD:1 M40:GATE 1.16601e-18 
c_1029 VDD:1 M39:GATE 3.56549e-18 
c_1030 VDD:1 M38:GATE 1.80066e-18 
c_1031 VDD:1 M41:GATE 5.38625e-19 
c_1032 VDD:1 M43:GATE 2.42927e-19 
c_1033 VDD:1 M42:GATE 1.16929e-18 
c_1034 VDD:1 0 2.74729e-17 
c_1035 VDD:2 M30:GATE 1.60854e-19 
c_1036 VDD:2 M31:GATE 1.22708e-19 
c_1037 VDD:2 M44:GATE 1.35814e-19 
c_1038 VDD:2 M46:GATE 1.30417e-19 
c_1039 VDD:2 M45:GATE 1.64815e-19 
c_1040 VDD:2 M36:SRC 6.266e-20 
c_1041 VDD:2 M34:GATE 6.52082e-20 
c_1042 VDD:2 M57:GATE 9.8175e-19 
c_1043 VDD:2 SDN:1 1.63347e-19 
c_1044 VDD:2 M58:GATE 1.67269e-18 
c_1045 VDD:2 N_56:1 1.45979e-18 
c_1046 VDD:2 N_15:3 8.83875e-17 
c_1047 VDD:2 SDN 5.44577e-19 
c_1048 VDD:2 N_15:1 6.8301e-19 
c_1049 VDD:2 M52:DRN 8.78699e-18 
c_1050 VDD:2 Q 4.08412e-17 
c_1051 VDD:2 M6:DRN 1.29566e-19 
c_1052 VDD:2 M50:DRN 7.36381e-19 
c_1053 VDD:2 M54:GATE 1.25816e-18 
c_1054 VDD:2 M53:GATE 1.10233e-18 
c_1055 VDD:2 M33:GATE 1.8851e-18 
c_1056 VDD:2 M37:GATE 4.4488e-19 
c_1057 VDD:2 M40:GATE 1.84766e-19 
c_1058 VDD:2 M39:GATE 9.03123e-20 
c_1059 VDD:2 M38:GATE 6.47945e-19 
c_1060 VDD:2 M56:GATE 2.47113e-18 
c_1061 VDD:2 M55:GATE 1.72217e-18 
c_1062 VDD:2 M52:GATE 9.96779e-19 
c_1063 VDD:2 M51:GATE 8.38278e-19 
c_1064 VDD:2 M50:GATE 1.14513e-18 
c_1065 VDD:2 M49:GATE 7.42903e-18 
c_1066 VDD:2 M43:GATE 1.9583e-18 
c_1067 VDD:2 0 1.89788e-17 
c_1068 VDD:3 M30:DRN 3.24711e-19 
c_1069 VDD:3 M20:DRN 8.26434e-21 
c_1070 VDD:3 M46:GATE 2.737e-20 
c_1071 VDD:3 M45:GATE 5.20462e-17 
c_1072 VDD:3 N_73:1 6.0819e-20 
c_1073 VDD:3 M34:GATE 7.02039e-19 
c_1074 VDD:3 M35:GATE 7.0165e-19 
c_1075 VDD:3 M57:GATE 4.45671e-19 
c_1076 VDD:3 SDN:1 8.33879e-20 
c_1077 VDD:3 M58:GATE 2.70832e-19 
c_1078 VDD:3 N_56:1 7.46934e-21 
c_1079 VDD:3 M54:GATE 2.05379e-19 
c_1080 VDD:3 M53:GATE 2.54759e-19 
c_1081 VDD:3 M56:GATE 5.10972e-19 
c_1082 VDD:3 M55:GATE 6.02877e-19 
c_1083 VDD:3 M52:GATE 2.05379e-19 
c_1084 VDD:3 M51:GATE 2.54759e-19 
c_1085 VDD:3 M50:GATE 2.05379e-19 
c_1086 VDD:3 M49:GATE 2.54759e-19 
c_1087 VDD:3 M43:GATE 9.18284e-19 
c_1088 VDD:3 0 2.23971e-17 
c_1089 M58:BULK M30:DRN 2.76231e-18 
c_1090 M58:BULK M25:GATE 2.6595e-18 
c_1091 M58:BULK M24:GATE 9.16553e-18 
c_1092 M58:BULK M24:SRC 4.3938e-19 
c_1093 M58:BULK D 1.61249e-19 
c_1094 M58:BULK M20:GATE 3.0385e-18 
c_1095 M58:BULK M30:GATE 3.72041e-17 
c_1096 M58:BULK SE 3.11589e-18 
c_1097 M58:BULK SI 3.05368e-18 
c_1098 M58:BULK M31:GATE 6.85003e-18 
c_1099 M58:BULK M44:GATE 5.25918e-18 
c_1100 M58:BULK M48:DRN 2.69957e-18 
c_1101 M58:BULK M48:SRC 1.84836e-18 
c_1102 M58:BULK M47:GATE 5.48442e-18 
c_1103 M58:BULK M45:GATE 1.8358e-17 
c_1104 M58:BULK M48:GATE 6.22318e-18 
c_1105 M58:BULK N_73:1 1.72724e-17 
c_1106 M58:BULK N_13:3 1.25064e-18 
c_1107 M58:BULK M9:GATE 4.65442e-19 
c_1108 M58:BULK M36:DRN 5.28031e-18 
c_1109 M58:BULK M34:GATE 1.27325e-17 
c_1110 M58:BULK M35:GATE 4.08164e-18 
c_1111 M58:BULK M35:DRN 5.82137e-18 
c_1112 M58:BULK N_62:1 7.83953e-18 
c_1113 M58:BULK M57:DRN 1.01976e-18 
c_1114 M58:BULK M57:GATE 1.98731e-17 
c_1115 M58:BULK SDN:1 3.56571e-17 
c_1116 M58:BULK M58:GATE 8.39268e-18 
c_1117 M58:BULK M58:SRC 1.87323e-18 
c_1118 M58:BULK M32:SRC 3.33718e-18 
c_1119 M58:BULK N_56:1 1.98783e-17 
c_1120 M58:BULK N_15:3 9.98471e-18 
c_1121 M58:BULK M15:SRC 7.59956e-19 
c_1122 M58:BULK CDN:1 1.74728e-18 
c_1123 M58:BULK M39:DRN 1.76868e-19 
c_1124 M58:BULK M43:DRN 4.11196e-19 
c_1125 M58:BULK SDN 4.82753e-18 
c_1126 M58:BULK N_13:1 3.3311e-18 
c_1127 M58:BULK N_13:2 3.53437e-18 
c_1128 M58:BULK N_15:1 1.50077e-18 
c_1129 M58:BULK M52:DRN 3.17687e-18 
c_1130 M58:BULK N_15:2 2.58692e-18 
c_1131 M58:BULK Q 7.71631e-18 
c_1132 M58:BULK M50:DRN 2.98131e-18 
c_1133 M58:BULK M54:GATE 5.53177e-18 
c_1134 M58:BULK M53:GATE 5.48294e-18 
c_1135 M58:BULK M33:GATE 2.77519e-18 
c_1136 M58:BULK M37:GATE 2.85509e-17 
c_1137 M58:BULK M27:GATE 2.83691e-18 
c_1138 M58:BULK M40:GATE 1.79845e-18 
c_1139 M58:BULK M39:GATE 1.21985e-18 
c_1140 M58:BULK M38:GATE 3.62492e-18 
c_1141 M58:BULK M56:GATE 4.3717e-18 
c_1142 M58:BULK M55:GATE 5.3583e-18 
c_1143 M58:BULK M52:GATE 3.18714e-18 
c_1144 M58:BULK M51:GATE 5.19817e-18 
c_1145 M58:BULK M50:GATE 5.10436e-18 
c_1146 M58:BULK M49:GATE 8.99524e-18 
c_1147 M58:BULK M41:GATE 3.5131e-18 
c_1148 M58:BULK CDN 1.2358e-18 
c_1149 M58:BULK M43:GATE 4.07421e-18 
c_1150 M58:BULK 0 1.27968e-17 
c_1151 VDD M30:DRN 1.17707e-18 
c_1152 VDD M24:SRC 1.87155e-18 
c_1153 VDD D 1.19852e-18 
c_1154 VDD M23:DRN 5.10407e-17 
c_1155 VDD M30:GATE 4.15036e-17 
c_1156 VDD SE 1.86409e-17 
c_1157 VDD SI 2.97787e-17 
c_1158 VDD M31:GATE 7.19413e-18 
c_1159 VDD M20:DRN 4.17651e-18 
c_1160 VDD M44:GATE 4.12737e-18 
c_1161 VDD M48:DRN 1.44101e-18 
c_1162 VDD M48:SRC 1.21912e-18 
c_1163 VDD M47:GATE 7.65814e-18 
c_1164 VDD M46:DRN 1.47146e-18 
c_1165 VDD M46:GATE 4.02137e-18 
c_1166 VDD M45:GATE 3.10254e-17 
c_1167 VDD M48:GATE 4.48048e-18 
c_1168 VDD N_73:1 2.08801e-16 
c_1169 VDD M28:SRC 2.77467e-18 
c_1170 VDD M36:SRC 2.7218e-19 
c_1171 VDD M36:DRN 3.64671e-19 
c_1172 VDD M34:GATE 5.69337e-19 
c_1173 VDD M57:DRN 1.86021e-20 
c_1174 VDD M57:GATE 4.22237e-18 
c_1175 VDD SDN:1 8.84785e-17 
c_1176 VDD M58:GATE 3.32672e-18 
c_1177 VDD M32:DRN 1.22128e-19 
c_1178 VDD N_56:1 1.76346e-17 
c_1179 VDD N_15:3 1.27182e-16 
c_1180 VDD M41:DRN 1.87387e-18 
c_1181 VDD M39:DRN 1.87387e-18 
c_1182 VDD SDN 1.92362e-19 
c_1183 VDD N_13:1 1.15541e-19 
c_1184 VDD N_15:1 6.05007e-19 
c_1185 VDD M52:DRN 2.80993e-18 
c_1186 VDD Q 8.72826e-17 
c_1187 VDD M50:DRN 2.80993e-18 
c_1188 VDD M54:GATE 7.23625e-18 
c_1189 VDD M53:GATE 7.56397e-18 
c_1190 VDD M33:GATE 2.06909e-16 
c_1191 VDD M40:GATE 1.90877e-18 
c_1192 VDD M39:GATE 5.2343e-19 
c_1193 VDD M38:GATE 6.23745e-19 
c_1194 VDD M56:GATE 6.9301e-18 
c_1195 VDD M55:GATE 6.92366e-18 
c_1196 VDD M52:GATE 7.07947e-18 
c_1197 VDD M51:GATE 6.84436e-18 
c_1198 VDD M50:GATE 6.86405e-18 
c_1199 VDD M49:GATE 6.561e-18 
c_1200 VDD M41:GATE 1.25717e-18 
c_1201 VDD M43:GATE 3.3907e-18 
c_1202 VDD M42:GATE 3.53601e-19 
c_1203 VDD 0 3.03908e-16 
c_1204 M55:DRN N_13:2 1.02597e-17 
c_1205 M55:DRN N_15:3 2.34327e-18 
c_1206 M55:DRN M56:GATE 8.3293e-19 
c_1207 M55:DRN M55:GATE 1.00916e-17 
c_1208 M55:DRN M54:GATE 1.00916e-17 
c_1209 M55:DRN M53:GATE 8.3293e-19 
c_1210 M55:DRN SDN:1 8.77326e-20 
c_1211 M55:DRN 0 6.5273e-18 
c_1212 M53:DRN Q 9.6272e-20 
c_1213 M53:DRN N_15:3 7.56232e-18 
c_1214 M53:DRN M54:GATE 8.3293e-19 
c_1215 M53:DRN M53:GATE 1.00916e-17 
c_1216 M53:DRN M52:GATE 1.00916e-17 
c_1217 M53:DRN M51:GATE 8.3293e-19 
c_1218 M53:DRN 0 3.70936e-18 
c_1219 M51:DRN Q 1.03274e-17 
c_1220 M51:DRN N_15:1 1.02252e-17 
c_1221 M51:DRN M52:GATE 8.3293e-19 
c_1222 M51:DRN M51:GATE 1.00916e-17 
c_1223 M51:DRN M50:GATE 1.002e-17 
c_1224 M51:DRN M49:GATE 1.12569e-18 
c_1225 M51:DRN 0 2.56554e-18 
c_1226 M56:SRC N_73:1 2.10147e-19 
c_1227 M56:SRC M57:GATE 1.06049e-22 
c_1228 M56:SRC SDN:1 2.28879e-17 
c_1229 M56:SRC M58:GATE 6.06794e-22 
c_1230 M56:SRC N_15:3 7.17862e-18 
c_1231 M56:SRC M18:SRC 9.72556e-19 
c_1232 M56:SRC N_13:1 8.02866e-18 
c_1233 M56:SRC M38:GATE 1.35909e-18 
c_1234 M56:SRC M56:GATE 2.17346e-17 
c_1235 M56:SRC M55:GATE 1.00502e-18 
c_1236 M56:SRC M43:GATE 1.13373e-17 
c_1237 M56:SRC 0 4.19952e-18 
c_1238 M49:DRN M49:GATE 3.4325e-17 
c_1239 M49:DRN M50:DRN 1.75167e-18 
c_1240 M49:DRN Q 1.38719e-18 
c_1241 M49:DRN M50:GATE 3.2182e-20 
c_1242 M49:DRN N_73:1 1.79599e-19 
c_1243 M49:DRN M6:DRN 8.04549e-20 
c_1244 M49:DRN 0 7.23538e-18 
c_1245 M57:SRC CDN:2 2.02488e-19 
c_1246 M57:SRC M3:DRN 1.14194e-19 
c_1247 M57:SRC M45:GATE 2.90962e-20 
c_1248 M57:SRC M36:DRN 2.21443e-22 
c_1249 M57:SRC M35:DRN 2.17028e-20 
c_1250 M57:SRC N_62:1 2.21278e-18 
c_1251 M57:SRC M57:GATE 1.34639e-17 
c_1252 M57:SRC M3:SRC 3.17548e-19 
c_1253 M57:SRC SDN:1 1.74207e-16 
c_1254 M57:SRC M58:GATE 1.4273e-17 
c_1255 M57:SRC M58:SRC 1.55028e-20 
c_1256 M57:SRC M2:DRN 3.41291e-19 
c_1257 M57:SRC M1:DRN 1.50365e-24 
c_1258 M57:SRC M32:SRC 4.02207e-20 
c_1259 M57:SRC M32:DRN 1.4283e-20 
c_1260 M57:SRC N_56:1 2.16217e-19 
c_1261 M57:SRC N_15:3 4.52232e-18 
c_1262 M57:SRC M41:DRN 1.9522e-20 
c_1263 M57:SRC CDN:1 5.98095e-21 
c_1264 M57:SRC M39:DRN 1.9522e-20 
c_1265 M57:SRC M18:SRC 1.48152e-19 
c_1266 M57:SRC M43:DRN 1.44071e-20 
c_1267 M57:SRC SDN 7.82941e-23 
c_1268 M57:SRC N_13:2 3.14971e-19 
c_1269 M57:SRC N_15:1 2.77371e-19 
c_1270 M57:SRC M52:DRN 1.07984e-18 
c_1271 M57:SRC Q 2.68015e-18 
c_1272 M57:SRC M50:DRN 1.07984e-18 
c_1273 M57:SRC M54:GATE 5.14431e-18 
c_1274 M57:SRC M53:GATE 3.77249e-18 
c_1275 M57:SRC M37:GATE 4.33618e-18 
c_1276 M57:SRC M40:GATE 1.70646e-19 
c_1277 M57:SRC M39:GATE 1.64958e-19 
c_1278 M57:SRC M38:GATE 1.70646e-19 
c_1279 M57:SRC M56:GATE 5.14333e-18 
c_1280 M57:SRC M55:GATE 5.14431e-18 
c_1281 M57:SRC M52:GATE 3.77154e-18 
c_1282 M57:SRC M51:GATE 5.14115e-18 
c_1283 M57:SRC M50:GATE 5.14115e-18 
c_1284 M57:SRC M49:GATE 5.13999e-18 
c_1285 M57:SRC M41:GATE 1.14199e-19 
c_1286 M57:SRC M43:GATE 7.23487e-20 
c_1287 M57:SRC M42:GATE 8.37457e-20 
c_1288 M57:SRC 0 3.19409e-17 
c_1289 M38:SRC N_73:1 3.08769e-19 
c_1290 M38:SRC SDN:1 2.13791e-17 
c_1291 M38:SRC M58:GATE 3.90949e-23 
c_1292 M38:SRC M58:SRC 6.71558e-23 
c_1293 M38:SRC N_15:3 2.48201e-17 
c_1294 M38:SRC M40:GATE 1.27185e-18 
c_1295 M38:SRC M39:GATE 1.50411e-17 
c_1296 M38:SRC M38:GATE 1.48393e-17 
c_1297 M38:SRC M43:GATE 2.92215e-18 
c_1298 M38:SRC 0 5.53644e-18 
c_1299 M42:SRC CDN:2 2.90582e-20 
c_1300 M42:SRC M36:SRC 2.30754e-20 
c_1301 M42:SRC M36:DRN 3.19515e-20 
c_1302 M42:SRC M57:GATE 1.06267e-20 
c_1303 M42:SRC SDN:1 6.59082e-17 
c_1304 M42:SRC M58:GATE 5.05821e-19 
c_1305 M42:SRC M58:SRC 1.38901e-19 
c_1306 M42:SRC M32:SRC 8.34889e-19 
c_1307 M42:SRC M32:DRN 1.44021e-17 
c_1308 M42:SRC N_56:1 9.94545e-18 
c_1309 M42:SRC M15:SRC 2.8177e-19 
c_1310 M42:SRC M41:DRN 5.69764e-18 
c_1311 M42:SRC M16:SRC 2.8009e-20 
c_1312 M42:SRC CDN:1 2.29397e-19 
c_1313 M42:SRC M39:DRN 2.55985e-21 
c_1314 M42:SRC N_13:1 1.916e-19 
c_1315 M42:SRC M37:GATE 3.53217e-18 
c_1316 M42:SRC M40:GATE 1.23654e-17 
c_1317 M42:SRC M39:GATE 1.2018e-18 
c_1318 M42:SRC M41:GATE 1.28882e-17 
c_1319 M42:SRC M43:GATE 4.39139e-20 
c_1320 M42:SRC M42:GATE 2.96083e-17 
c_1321 M42:SRC 0 1.15678e-17 
c_1322 M40:SRC SDN:1 1.82168e-18 
c_1323 M40:SRC M58:SRC 1.56396e-22 
c_1324 M40:SRC M32:SRC 8.13874e-23 
c_1325 M40:SRC N_56:1 2.067e-18 
c_1326 M40:SRC N_15:3 2.756e-18 
c_1327 M40:SRC M15:GATE 1.30604e-18 
c_1328 M40:SRC M16:SRC 2.92301e-18 
c_1329 M40:SRC CDN:1 1.97879e-19 
c_1330 M40:SRC M41:GATE 6.36711e-18 
c_1331 M40:SRC CDN 6.61723e-18 
c_1332 M40:SRC M42:GATE 7.29948e-19 
c_1333 M35:SRC M30:GATE 1.06049e-22 
c_1334 M35:SRC M46:GATE 1.58368e-20 
c_1335 M35:SRC M28:SRC 1.57735e-19 
c_1336 M35:SRC M36:SRC 8.22646e-20 
c_1337 M35:SRC M36:DRN 1.02501e-19 
c_1338 M35:SRC M34:GATE 1.55441e-17 
c_1339 M35:SRC M27:DRN 1.50337e-18 
c_1340 M35:SRC M35:GATE 1.44951e-17 
c_1341 M35:SRC M35:DRN 3.24259e-18 
c_1342 M35:SRC N_62:1 1.47999e-18 
c_1343 M35:SRC M57:DRN 2.34089e-18 
c_1344 M35:SRC M57:GATE 2.2832e-18 
c_1345 M35:SRC SDN:1 4.58595e-19 
c_1346 M35:SRC M58:GATE 5.25291e-20 
c_1347 M35:SRC M33:GATE 1.05219e-17 
c_1348 M35:SRC M56:GATE 7.95366e-22 
c_1349 M35:SRC 0 8.62994e-19 
c_1350 M47:DRN M22:GATE 7.51825e-24 
c_1351 M47:DRN M30:DRN 7.06446e-18 
c_1352 M47:DRN M23:GATE 1.20292e-23 
c_1353 M47:DRN M24:SRC 8.72245e-19 
c_1354 M47:DRN D 1.10085e-17 
c_1355 M47:DRN CDN:2 2.70657e-23 
c_1356 M47:DRN M23:DRN 4.9945e-20 
c_1357 M47:DRN M44:DRN 3.00333e-18 
c_1358 M47:DRN M30:GATE 6.49047e-17 
c_1359 M47:DRN SE 8.41385e-23 
c_1360 M47:DRN SI 2.01552e-20 
c_1361 M47:DRN M31:GATE 1.80799e-18 
c_1362 M47:DRN M20:DRN 2.39294e-18 
c_1363 M47:DRN M3:DRN 4.61007e-20 
c_1364 M47:DRN M44:GATE 1.80752e-18 
c_1365 M47:DRN M48:DRN 7.81094e-18 
c_1366 M47:DRN M48:SRC 8.51738e-18 
c_1367 M47:DRN M47:GATE 2.53388e-17 
c_1368 M47:DRN CP 2.69607e-19 
c_1369 M47:DRN M46:DRN 4.73381e-17 
c_1370 M47:DRN M46:GATE 1.39152e-17 
c_1371 M47:DRN M45:GATE 4.76303e-17 
c_1372 M47:DRN M48:GATE 2.87253e-17 
c_1373 M47:DRN N_73:1 5.4059e-18 
c_1374 M47:DRN M28:SRC 4.74439e-19 
c_1375 M47:DRN M36:SRC 6.98696e-18 
c_1376 M47:DRN M36:DRN 2.63143e-18 
c_1377 M47:DRN M33:DRN 5.87012e-19 
c_1378 M47:DRN M34:DRN 4.02554e-18 
c_1379 M47:DRN M34:GATE 3.19634e-18 
c_1380 M47:DRN M35:GATE 1.52044e-19 
c_1381 M47:DRN M35:DRN 2.37161e-18 
c_1382 M47:DRN M57:DRN 6.95523e-18 
c_1383 M47:DRN M57:GATE 3.79219e-18 
c_1384 M47:DRN M3:SRC 2.22334e-19 
c_1385 M47:DRN SDN:1 1.17849e-16 
c_1386 M47:DRN M58:GATE 1.1579e-19 
c_1387 M47:DRN M58:SRC 4.49015e-18 
c_1388 M47:DRN M2:DRN 2.62583e-20 
c_1389 M47:DRN M2:SRC 3.44424e-20 
c_1390 M47:DRN M1:DRN 5.76453e-20 
c_1391 M47:DRN M32:SRC 1.23029e-18 
c_1392 M47:DRN M32:DRN 8.66206e-19 
c_1393 M47:DRN N_15:3 4.77685e-20 
c_1394 M47:DRN M41:DRN 8.6913e-20 
c_1395 M47:DRN M16:SRC 3.40963e-21 
c_1396 M47:DRN M39:DRN 3.51071e-18 
c_1397 M47:DRN M18:SRC 1.47734e-19 
c_1398 M47:DRN M43:DRN 3.22166e-18 
c_1399 M47:DRN N_13:2 1.24326e-19 
c_1400 M47:DRN N_15:1 1.24326e-19 
c_1401 M47:DRN M8:DRN 3.81007e-20 
c_1402 M47:DRN M52:DRN 1.02793e-17 
c_1403 M47:DRN M6:DRN 3.81007e-20 
c_1404 M47:DRN M50:DRN 1.02793e-17 
c_1405 M47:DRN M54:GATE 4.35799e-18 
c_1406 M47:DRN M53:GATE 5.29123e-18 
c_1407 M47:DRN M33:GATE 5.39641e-17 
c_1408 M47:DRN M27:GATE 4.65738e-23 
c_1409 M47:DRN M40:GATE 1.65019e-18 
c_1410 M47:DRN M39:GATE 1.64713e-18 
c_1411 M47:DRN M38:GATE 1.64713e-18 
c_1412 M47:DRN M56:GATE 4.35799e-18 
c_1413 M47:DRN M55:GATE 4.35799e-18 
c_1414 M47:DRN M52:GATE 5.29123e-18 
c_1415 M47:DRN M51:GATE 4.35799e-18 
c_1416 M47:DRN M50:GATE 4.35799e-18 
c_1417 M47:DRN M49:GATE 4.35799e-18 
c_1418 M47:DRN 0 2.98357e-16 
c_1419 M46:SRC M33:GATE 2.61964e-19 
c_1420 M46:SRC M36:SRC 5.20866e-20 
c_1421 M46:SRC N_73:1 3.10923e-18 
c_1422 M46:SRC M30:GATE 7.85103e-20 
c_1423 M46:SRC M46:GATE 8.49554e-18 
c_1424 M46:SRC M45:GATE 1.19815e-17 
c_1425 M46:SRC M20:DRN 3.38023e-18 
c_1426 M46:SRC 0 2.36727e-18 
c_1427 M31:DRN M30:DRN 1.04894e-18 
c_1428 M31:DRN M23:GATE 7.21752e-23 
c_1429 M31:DRN M23:DRN 5.77789e-19 
c_1430 M31:DRN M30:GATE 6.33618e-18 
c_1431 M31:DRN SE 2.27e-17 
c_1432 M31:DRN SI 9.92403e-19 
c_1433 M31:DRN M31:GATE 1.92692e-17 
c_1434 M31:DRN M44:GATE 1.08677e-18 
c_1435 M31:DRN M48:DRN 5.93543e-19 
c_1436 M31:DRN M48:SRC 2.28381e-21 
c_1437 M31:DRN 0 1.46525e-18 

.ENDS
